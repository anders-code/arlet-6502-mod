`ifdef TT_SYNTH
    `define USE_ASYNC_RESET 1
    `define NO_TIMESCALE 1
`endif
