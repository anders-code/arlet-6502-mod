module tt_um_anders_tt_6502 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire net126;
 wire clknet_0_clk;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire net104;
 wire \cpu_inst.ABH[0] ;
 wire \cpu_inst.ABH[1] ;
 wire \cpu_inst.ABH[2] ;
 wire \cpu_inst.ABH[3] ;
 wire \cpu_inst.ABH[4] ;
 wire \cpu_inst.ABH[5] ;
 wire \cpu_inst.ABH[6] ;
 wire \cpu_inst.ABH[7] ;
 wire \cpu_inst.ABL[0] ;
 wire \cpu_inst.ABL[1] ;
 wire \cpu_inst.ABL[2] ;
 wire \cpu_inst.ABL[3] ;
 wire \cpu_inst.ABL[4] ;
 wire \cpu_inst.ABL[5] ;
 wire \cpu_inst.ABL[6] ;
 wire \cpu_inst.ABL[7] ;
 wire \cpu_inst.ADD[0] ;
 wire \cpu_inst.ADD[1] ;
 wire \cpu_inst.ADD[2] ;
 wire \cpu_inst.ADD[3] ;
 wire \cpu_inst.ADD[4] ;
 wire \cpu_inst.ADD[5] ;
 wire \cpu_inst.ADD[6] ;
 wire \cpu_inst.ADD[7] ;
 wire \cpu_inst.ALU.AI7 ;
 wire \cpu_inst.ALU.BI7 ;
 wire \cpu_inst.ALU.CO ;
 wire \cpu_inst.ALU.HC ;
 wire \cpu_inst.AXYS[0][0] ;
 wire \cpu_inst.AXYS[0][1] ;
 wire \cpu_inst.AXYS[0][2] ;
 wire \cpu_inst.AXYS[0][3] ;
 wire \cpu_inst.AXYS[0][4] ;
 wire \cpu_inst.AXYS[0][5] ;
 wire \cpu_inst.AXYS[0][6] ;
 wire \cpu_inst.AXYS[0][7] ;
 wire \cpu_inst.AXYS[1][0] ;
 wire \cpu_inst.AXYS[1][1] ;
 wire \cpu_inst.AXYS[1][2] ;
 wire \cpu_inst.AXYS[1][3] ;
 wire \cpu_inst.AXYS[1][4] ;
 wire \cpu_inst.AXYS[1][5] ;
 wire \cpu_inst.AXYS[1][6] ;
 wire \cpu_inst.AXYS[1][7] ;
 wire \cpu_inst.AXYS[2][0] ;
 wire \cpu_inst.AXYS[2][1] ;
 wire \cpu_inst.AXYS[2][2] ;
 wire \cpu_inst.AXYS[2][3] ;
 wire \cpu_inst.AXYS[2][4] ;
 wire \cpu_inst.AXYS[2][5] ;
 wire \cpu_inst.AXYS[2][6] ;
 wire \cpu_inst.AXYS[2][7] ;
 wire \cpu_inst.AXYS[3][0] ;
 wire \cpu_inst.AXYS[3][1] ;
 wire \cpu_inst.AXYS[3][2] ;
 wire \cpu_inst.AXYS[3][3] ;
 wire \cpu_inst.AXYS[3][4] ;
 wire \cpu_inst.AXYS[3][5] ;
 wire \cpu_inst.AXYS[3][6] ;
 wire \cpu_inst.AXYS[3][7] ;
 wire \cpu_inst.C ;
 wire \cpu_inst.D ;
 wire \cpu_inst.DI[0] ;
 wire \cpu_inst.DI[1] ;
 wire \cpu_inst.DI[2] ;
 wire \cpu_inst.DI[3] ;
 wire \cpu_inst.DI[4] ;
 wire \cpu_inst.DI[5] ;
 wire \cpu_inst.DI[6] ;
 wire \cpu_inst.DI[7] ;
 wire \cpu_inst.I ;
 wire \cpu_inst.IRHOLD[0] ;
 wire \cpu_inst.IRHOLD[1] ;
 wire \cpu_inst.IRHOLD[2] ;
 wire \cpu_inst.IRHOLD[3] ;
 wire \cpu_inst.IRHOLD[4] ;
 wire \cpu_inst.IRHOLD[5] ;
 wire \cpu_inst.IRHOLD[6] ;
 wire \cpu_inst.IRHOLD[7] ;
 wire \cpu_inst.IRHOLD_valid ;
 wire \cpu_inst.N ;
 wire \cpu_inst.NMI_1 ;
 wire \cpu_inst.NMI_edge ;
 wire \cpu_inst.PC[0] ;
 wire \cpu_inst.PC[10] ;
 wire \cpu_inst.PC[11] ;
 wire \cpu_inst.PC[12] ;
 wire \cpu_inst.PC[13] ;
 wire \cpu_inst.PC[14] ;
 wire \cpu_inst.PC[15] ;
 wire \cpu_inst.PC[1] ;
 wire \cpu_inst.PC[2] ;
 wire \cpu_inst.PC[3] ;
 wire \cpu_inst.PC[4] ;
 wire \cpu_inst.PC[5] ;
 wire \cpu_inst.PC[6] ;
 wire \cpu_inst.PC[7] ;
 wire \cpu_inst.PC[8] ;
 wire \cpu_inst.PC[9] ;
 wire \cpu_inst.V ;
 wire \cpu_inst.Z ;
 wire \cpu_inst.adc_bcd ;
 wire \cpu_inst.adc_sbc ;
 wire \cpu_inst.adj_bcd ;
 wire \cpu_inst.backwards ;
 wire \cpu_inst.bit_ins ;
 wire \cpu_inst.clc ;
 wire \cpu_inst.cld ;
 wire \cpu_inst.cli ;
 wire \cpu_inst.clv ;
 wire \cpu_inst.compare ;
 wire \cpu_inst.cond_code[0] ;
 wire \cpu_inst.cond_code[1] ;
 wire \cpu_inst.cond_code[2] ;
 wire \cpu_inst.dst_reg[0] ;
 wire \cpu_inst.dst_reg[1] ;
 wire \cpu_inst.inc ;
 wire \cpu_inst.index_y ;
 wire \cpu_inst.load_only ;
 wire \cpu_inst.load_reg ;
 wire \cpu_inst.op[0] ;
 wire \cpu_inst.op[1] ;
 wire \cpu_inst.op[2] ;
 wire \cpu_inst.op[3] ;
 wire \cpu_inst.php ;
 wire \cpu_inst.plp ;
 wire \cpu_inst.res ;
 wire \cpu_inst.rotate ;
 wire \cpu_inst.sec ;
 wire \cpu_inst.sed ;
 wire \cpu_inst.sei ;
 wire \cpu_inst.shift ;
 wire \cpu_inst.shift_right ;
 wire \cpu_inst.src_reg[0] ;
 wire \cpu_inst.src_reg[1] ;
 wire \cpu_inst.state[0] ;
 wire \cpu_inst.state[1] ;
 wire \cpu_inst.state[2] ;
 wire \cpu_inst.state[3] ;
 wire \cpu_inst.state[4] ;
 wire \cpu_inst.state[5] ;
 wire \cpu_inst.store ;
 wire \cpu_inst.write_back ;
 wire \spi_sram_master_inst.counter[0] ;
 wire \spi_sram_master_inst.counter[1] ;
 wire \spi_sram_master_inst.counter[2] ;
 wire \spi_sram_master_inst.counter[3] ;
 wire \spi_sram_master_inst.counter[4] ;
 wire \spi_sram_master_inst.counter_done ;
 wire \spi_sram_master_inst.cs_n ;
 wire \spi_sram_master_inst.cs_n_sm ;
 wire \spi_sram_master_inst.data[10] ;
 wire \spi_sram_master_inst.data[11] ;
 wire \spi_sram_master_inst.data[12] ;
 wire \spi_sram_master_inst.data[13] ;
 wire \spi_sram_master_inst.data[14] ;
 wire \spi_sram_master_inst.data[15] ;
 wire \spi_sram_master_inst.data[16] ;
 wire \spi_sram_master_inst.data[17] ;
 wire \spi_sram_master_inst.data[18] ;
 wire \spi_sram_master_inst.data[19] ;
 wire \spi_sram_master_inst.data[20] ;
 wire \spi_sram_master_inst.data[21] ;
 wire \spi_sram_master_inst.data[22] ;
 wire \spi_sram_master_inst.data[23] ;
 wire \spi_sram_master_inst.data[24] ;
 wire \spi_sram_master_inst.data[25] ;
 wire \spi_sram_master_inst.data[26] ;
 wire \spi_sram_master_inst.data[27] ;
 wire \spi_sram_master_inst.data[28] ;
 wire \spi_sram_master_inst.data[29] ;
 wire \spi_sram_master_inst.data[30] ;
 wire \spi_sram_master_inst.data[31] ;
 wire \spi_sram_master_inst.data[32] ;
 wire \spi_sram_master_inst.data[33] ;
 wire \spi_sram_master_inst.data[34] ;
 wire \spi_sram_master_inst.data[35] ;
 wire \spi_sram_master_inst.data[36] ;
 wire \spi_sram_master_inst.data[37] ;
 wire \spi_sram_master_inst.data[38] ;
 wire \spi_sram_master_inst.data[39] ;
 wire \spi_sram_master_inst.data[8] ;
 wire \spi_sram_master_inst.data[9] ;
 wire \spi_sram_master_inst.dout ;
 wire \spi_sram_master_inst.state[0] ;
 wire \spi_sram_master_inst.state[1] ;
 wire \spi_sram_master_inst.state[2] ;
 wire \spi_sram_master_inst.state[3] ;
 wire \spi_sram_master_inst.state[4] ;
 wire \spi_sram_master_inst.state[5] ;
 wire \spi_sram_master_inst.state[6] ;
 wire \spi_sram_master_inst.state[7] ;
 wire net123;
 wire net124;
 wire net105;
 wire net125;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;

 sky130_fd_sc_hd__inv_2 _1062_ (.A(\cpu_inst.NMI_edge ),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(net85),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(net81),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(\cpu_inst.AXYS[2][0] ),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(\cpu_inst.AXYS[3][0] ),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(\cpu_inst.C ),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(\cpu_inst.clc ),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(net207),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(\cpu_inst.cld ),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(\cpu_inst.php ),
    .Y(_0508_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(net205),
    .Y(_0509_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(net245),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_2 _2123__2 (.A(clknet_4_5_0_clk),
    .Y(net126));
 sky130_fd_sc_hd__a21o_1 _1075_ (.A1(net209),
    .A2(_0506_),
    .B1(\spi_sram_master_inst.state[2] ),
    .X(_0005_));
 sky130_fd_sc_hd__nor2_2 _1076_ (.A(\spi_sram_master_inst.state[0] ),
    .B(net232),
    .Y(_0511_));
 sky130_fd_sc_hd__a21bo_1 _1077_ (.A1(net223),
    .A2(_0506_),
    .B1_N(_0511_),
    .X(_0004_));
 sky130_fd_sc_hd__or4_1 _1078_ (.A(\spi_sram_master_inst.state[5] ),
    .B(\spi_sram_master_inst.state[0] ),
    .C(\spi_sram_master_inst.state[7] ),
    .D(\spi_sram_master_inst.state[3] ),
    .X(\spi_sram_master_inst.cs_n_sm ));
 sky130_fd_sc_hd__or2_1 _1079_ (.A(\spi_sram_master_inst.counter[0] ),
    .B(\spi_sram_master_inst.counter[1] ),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _1080_ (.A(\spi_sram_master_inst.counter[2] ),
    .B(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__a21oi_1 _1081_ (.A1(\spi_sram_master_inst.counter[2] ),
    .A2(_0512_),
    .B1(\spi_sram_master_inst.state[2] ),
    .Y(_0514_));
 sky130_fd_sc_hd__a21o_1 _1082_ (.A1(_0513_),
    .A2(_0514_),
    .B1(\spi_sram_master_inst.state[1] ),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _1083_ (.A(_0511_),
    .B(_0515_),
    .Y(_0006_));
 sky130_fd_sc_hd__or2_1 _1084_ (.A(\spi_sram_master_inst.counter[3] ),
    .B(_0513_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_1 _1085_ (.A(\spi_sram_master_inst.counter[3] ),
    .B(_0513_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_1 _1086_ (.A(\spi_sram_master_inst.state[1] ),
    .B(\spi_sram_master_inst.state[2] ),
    .Y(_0518_));
 sky130_fd_sc_hd__a21bo_1 _1087_ (.A1(_0516_),
    .A2(_0517_),
    .B1_N(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__nand2_1 _1088_ (.A(_0511_),
    .B(_0519_),
    .Y(_0007_));
 sky130_fd_sc_hd__and3_1 _1089_ (.A(\spi_sram_master_inst.counter[4] ),
    .B(_0516_),
    .C(_0518_),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_1 _1090_ (.A(_0511_),
    .B(_0518_),
    .Y(_0521_));
 sky130_fd_sc_hd__nor3_1 _1091_ (.A(net130),
    .B(_0516_),
    .C(_0521_),
    .Y(_0187_));
 sky130_fd_sc_hd__or3b_1 _1092_ (.A(_0520_),
    .B(_0187_),
    .C_N(_0511_),
    .X(_0008_));
 sky130_fd_sc_hd__nor2_2 _1093_ (.A(\spi_sram_master_inst.state[5] ),
    .B(\spi_sram_master_inst.state[0] ),
    .Y(_0522_));
 sky130_fd_sc_hd__or2_1 _1094_ (.A(\spi_sram_master_inst.state[5] ),
    .B(\spi_sram_master_inst.state[0] ),
    .X(_0523_));
 sky130_fd_sc_hd__and2b_1 _1095_ (.A_N(net86),
    .B(net85),
    .X(_0524_));
 sky130_fd_sc_hd__nand2b_1 _1096_ (.A_N(\cpu_inst.state[4] ),
    .B(net85),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_1 _1097_ (.A(net87),
    .B(net90),
    .Y(_0526_));
 sky130_fd_sc_hd__nand4_2 _1098_ (.A(net94),
    .B(net92),
    .C(net88),
    .D(net90),
    .Y(_0527_));
 sky130_fd_sc_hd__nor2_1 _1099_ (.A(net54),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_1 _1100_ (.A(\cpu_inst.NMI_edge ),
    .B(net2),
    .Y(_0529_));
 sky130_fd_sc_hd__a21o_2 _1101_ (.A1(_0499_),
    .A2(\cpu_inst.I ),
    .B1(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_4 _1102_ (.A0(net98),
    .A1(\cpu_inst.IRHOLD[2] ),
    .S(net75),
    .X(_0531_));
 sky130_fd_sc_hd__nand2_1 _1103_ (.A(net49),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__mux2_2 _1104_ (.A0(net97),
    .A1(\cpu_inst.IRHOLD[3] ),
    .S(net75),
    .X(_0533_));
 sky130_fd_sc_hd__nor2_1 _1105_ (.A(_0532_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__nor2_1 _1106_ (.A(net86),
    .B(net85),
    .Y(_0535_));
 sky130_fd_sc_hd__or2_1 _1107_ (.A(net86),
    .B(net85),
    .X(_0536_));
 sky130_fd_sc_hd__or4bb_4 _1108_ (.A(net94),
    .B(net92),
    .C_N(net87),
    .D_N(net89),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_1 _1109_ (.A(net69),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__nor2_2 _1110_ (.A(net52),
    .B(_0537_),
    .Y(_0539_));
 sky130_fd_sc_hd__or2_2 _1111_ (.A(net52),
    .B(_0537_),
    .X(_0540_));
 sky130_fd_sc_hd__nor2_1 _1112_ (.A(net71),
    .B(net47),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _1113_ (.A(net57),
    .B(net48),
    .Y(_0542_));
 sky130_fd_sc_hd__mux2_2 _1114_ (.A0(\cpu_inst.DI[4] ),
    .A1(\cpu_inst.IRHOLD[4] ),
    .S(net75),
    .X(_0543_));
 sky130_fd_sc_hd__inv_2 _1115_ (.A(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__and2_2 _1116_ (.A(net49),
    .B(_0543_),
    .X(_0545_));
 sky130_fd_sc_hd__nand2_2 _1117_ (.A(net49),
    .B(_0543_),
    .Y(_0546_));
 sky130_fd_sc_hd__a32o_1 _1118_ (.A1(_0534_),
    .A2(net30),
    .A3(_0546_),
    .B1(_0528_),
    .B2(net68),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_2 _1119_ (.A(_0527_),
    .B(net52),
    .Y(_0548_));
 sky130_fd_sc_hd__nand4b_2 _1120_ (.A_N(net93),
    .B(net92),
    .C(net87),
    .D(net90),
    .Y(_0549_));
 sky130_fd_sc_hd__nor2_1 _1121_ (.A(net52),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__mux2_1 _1122_ (.A0(_0548_),
    .A1(_0550_),
    .S(net57),
    .X(_0551_));
 sky130_fd_sc_hd__or2_1 _1123_ (.A(_0547_),
    .B(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__nand4b_4 _1124_ (.A_N(net88),
    .B(net89),
    .C(net93),
    .D(net91),
    .Y(_0553_));
 sky130_fd_sc_hd__nor2_4 _1125_ (.A(net55),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__or2_2 _1126_ (.A(net55),
    .B(_0553_),
    .X(_0555_));
 sky130_fd_sc_hd__or4bb_4 _1127_ (.A(net93),
    .B(net88),
    .C_N(net89),
    .D_N(net91),
    .X(_0556_));
 sky130_fd_sc_hd__or2_1 _1128_ (.A(net55),
    .B(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__inv_2 _1129_ (.A(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__mux2_1 _1130_ (.A0(_0555_),
    .A1(_0557_),
    .S(net61),
    .X(_0559_));
 sky130_fd_sc_hd__nand2b_1 _1131_ (.A_N(net85),
    .B(net86),
    .Y(_0560_));
 sky130_fd_sc_hd__or2_1 _1132_ (.A(net70),
    .B(net50),
    .X(_0561_));
 sky130_fd_sc_hd__or2_2 _1133_ (.A(net58),
    .B(net50),
    .X(_0562_));
 sky130_fd_sc_hd__o22ai_1 _1134_ (.A1(_0556_),
    .A2(_0561_),
    .B1(_0562_),
    .B2(_0553_),
    .Y(_0563_));
 sky130_fd_sc_hd__or3b_1 _1135_ (.A(_0552_),
    .B(_0563_),
    .C_N(_0559_),
    .X(_0564_));
 sky130_fd_sc_hd__or4bb_4 _1136_ (.A(net93),
    .B(net89),
    .C_N(net88),
    .D_N(net91),
    .X(_0565_));
 sky130_fd_sc_hd__nor2_2 _1137_ (.A(net53),
    .B(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__and4b_2 _1138_ (.A_N(net89),
    .B(net88),
    .C(net91),
    .D(net93),
    .X(_0567_));
 sky130_fd_sc_hd__and2_2 _1139_ (.A(_0535_),
    .B(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_1 _1140_ (.A(_0535_),
    .B(_0567_),
    .Y(_0569_));
 sky130_fd_sc_hd__mux2_1 _1141_ (.A0(net46),
    .A1(_0568_),
    .S(net70),
    .X(_0570_));
 sky130_fd_sc_hd__or2_2 _1142_ (.A(net51),
    .B(_0565_),
    .X(_0571_));
 sky130_fd_sc_hd__nand2b_4 _1143_ (.A_N(net50),
    .B(_0567_),
    .Y(_0572_));
 sky130_fd_sc_hd__o22ai_1 _1144_ (.A1(_0561_),
    .A2(_0565_),
    .B1(_0572_),
    .B2(net58),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_2 _1145_ (.A(_0524_),
    .B(_0567_),
    .Y(_0574_));
 sky130_fd_sc_hd__or2_2 _1146_ (.A(net55),
    .B(_0565_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _1147_ (.A0(_0574_),
    .A1(_0575_),
    .S(net56),
    .X(_0576_));
 sky130_fd_sc_hd__or3b_1 _1148_ (.A(_0570_),
    .B(_0573_),
    .C_N(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_2 _1149_ (.A(net52),
    .B(_0553_),
    .Y(_0578_));
 sky130_fd_sc_hd__nor2_1 _1150_ (.A(_0549_),
    .B(net50),
    .Y(_0579_));
 sky130_fd_sc_hd__nor2_1 _1151_ (.A(_0527_),
    .B(net50),
    .Y(_0580_));
 sky130_fd_sc_hd__mux2_1 _1152_ (.A0(_0579_),
    .A1(_0580_),
    .S(net68),
    .X(_0581_));
 sky130_fd_sc_hd__nor2_1 _1153_ (.A(net53),
    .B(_0556_),
    .Y(_0582_));
 sky130_fd_sc_hd__xor2_2 _1154_ (.A(\cpu_inst.backwards ),
    .B(net84),
    .X(_0583_));
 sky130_fd_sc_hd__and3_1 _1155_ (.A(net57),
    .B(net42),
    .C(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__a211o_1 _1156_ (.A1(net69),
    .A2(net43),
    .B1(_0581_),
    .C1(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__or4b_4 _1157_ (.A(net93),
    .B(net87),
    .C(net90),
    .D_N(net91),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _1158_ (.A(net52),
    .B(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__inv_2 _1159_ (.A(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__or4bb_4 _1160_ (.A(net88),
    .B(net89),
    .C_N(net93),
    .D_N(net91),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _1161_ (.A(net51),
    .B(_0586_),
    .Y(_0590_));
 sky130_fd_sc_hd__nor2_1 _1162_ (.A(net51),
    .B(_0589_),
    .Y(_0591_));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(_0590_),
    .A1(_0591_),
    .S(net71),
    .X(_0592_));
 sky130_fd_sc_hd__nor2_1 _1164_ (.A(net53),
    .B(_0589_),
    .Y(_0593_));
 sky130_fd_sc_hd__mux2_1 _1165_ (.A0(_0588_),
    .A1(_0593_),
    .S(net68),
    .X(_0594_));
 sky130_fd_sc_hd__or4b_4 _1166_ (.A(net93),
    .B(net91),
    .C(net88),
    .D_N(net89),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _1167_ (.A(net52),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_1 _1168_ (.A(_0528_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2b_1 _1170_ (.A_N(net92),
    .B(net94),
    .Y(_0599_));
 sky130_fd_sc_hd__or3_2 _1171_ (.A(net87),
    .B(net90),
    .C(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_2 _1172_ (.A(net55),
    .B(net51),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_2 _1173_ (.A(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__o21ai_1 _1174_ (.A1(_0600_),
    .A2(_0601_),
    .B1(_0597_),
    .Y(_0603_));
 sky130_fd_sc_hd__nor2_1 _1175_ (.A(net54),
    .B(_0589_),
    .Y(_0604_));
 sky130_fd_sc_hd__and2_1 _1176_ (.A(net68),
    .B(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__a31o_1 _1177_ (.A1(\cpu_inst.write_back ),
    .A2(net57),
    .A3(_0603_),
    .B1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__or4_1 _1178_ (.A(_0585_),
    .B(_0592_),
    .C(_0594_),
    .D(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__or3_1 _1179_ (.A(_0564_),
    .B(_0577_),
    .C(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__nor2_1 _1180_ (.A(_0526_),
    .B(_0599_),
    .Y(_0609_));
 sky130_fd_sc_hd__a21o_1 _1181_ (.A1(net69),
    .A2(_0609_),
    .B1(_0538_),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_1 _1182_ (.A(net49),
    .B(_0533_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _1183_ (.A(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__or2_2 _1184_ (.A(_0531_),
    .B(_0611_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_2 _1185_ (.A0(net100),
    .A1(\cpu_inst.IRHOLD[0] ),
    .S(net75),
    .X(_0614_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(net49),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__mux2_2 _1187_ (.A0(net99),
    .A1(\cpu_inst.IRHOLD[1] ),
    .S(net75),
    .X(_0616_));
 sky130_fd_sc_hd__or2_2 _1188_ (.A(_0615_),
    .B(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _1189_ (.A(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _1190_ (.A(_0611_),
    .B(_0615_),
    .Y(_0619_));
 sky130_fd_sc_hd__mux2_2 _1191_ (.A0(net95),
    .A1(\cpu_inst.IRHOLD[7] ),
    .S(net75),
    .X(_0620_));
 sky130_fd_sc_hd__and2_1 _1192_ (.A(net49),
    .B(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__nand2_4 _1193_ (.A(_0530_),
    .B(_0620_),
    .Y(_0622_));
 sky130_fd_sc_hd__o32a_1 _1194_ (.A1(_0531_),
    .A2(_0619_),
    .A3(_0622_),
    .B1(_0613_),
    .B2(_0617_),
    .X(_0623_));
 sky130_fd_sc_hd__and3b_1 _1195_ (.A_N(_0623_),
    .B(net48),
    .C(_0546_),
    .X(_0624_));
 sky130_fd_sc_hd__nor2_1 _1196_ (.A(net50),
    .B(_0595_),
    .Y(_0625_));
 sky130_fd_sc_hd__or4_1 _1197_ (.A(net84),
    .B(\cpu_inst.store ),
    .C(net50),
    .D(_0595_),
    .X(_0626_));
 sky130_fd_sc_hd__or2_2 _1198_ (.A(_0593_),
    .B(_0625_),
    .X(_0627_));
 sky130_fd_sc_hd__nor3b_1 _1199_ (.A(net84),
    .B(\cpu_inst.store ),
    .C_N(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__o2bb2a_1 _1200_ (.A1_N(\cpu_inst.write_back ),
    .A2_N(_0626_),
    .B1(_0628_),
    .B2(_0603_),
    .X(_0629_));
 sky130_fd_sc_hd__and2_1 _1201_ (.A(_0601_),
    .B(_0609_),
    .X(_0630_));
 sky130_fd_sc_hd__nor3_2 _1202_ (.A(net87),
    .B(net50),
    .C(_0599_),
    .Y(_0631_));
 sky130_fd_sc_hd__nor2_1 _1203_ (.A(net54),
    .B(_0549_),
    .Y(_0632_));
 sky130_fd_sc_hd__or3_1 _1204_ (.A(\cpu_inst.state[4] ),
    .B(_0526_),
    .C(_0599_),
    .X(_0633_));
 sky130_fd_sc_hd__nor2_2 _1205_ (.A(net85),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(_0535_),
    .B(_0609_),
    .Y(_0635_));
 sky130_fd_sc_hd__or3_1 _1207_ (.A(_0630_),
    .B(_0631_),
    .C(net38),
    .X(_0636_));
 sky130_fd_sc_hd__o31a_1 _1208_ (.A1(_0624_),
    .A2(_0629_),
    .A3(_0636_),
    .B1(net57),
    .X(_0637_));
 sky130_fd_sc_hd__a221o_1 _1209_ (.A1(_0601_),
    .A2(_0610_),
    .B1(_0634_),
    .B2(net69),
    .C1(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__or4bb_4 _1210_ (.A(net91),
    .B(net88),
    .C_N(net89),
    .D_N(net93),
    .X(_0639_));
 sky130_fd_sc_hd__nor2_1 _1211_ (.A(net55),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__or2_1 _1212_ (.A(net54),
    .B(_0639_),
    .X(_0641_));
 sky130_fd_sc_hd__nor2_1 _1213_ (.A(net59),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand2_2 _1214_ (.A(net49),
    .B(_0616_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_4 _1215_ (.A(_0615_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _1216_ (.A(_0532_),
    .B(_0611_),
    .Y(_0645_));
 sky130_fd_sc_hd__nor2_1 _1217_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _1218_ (.A(net30),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__mux2_1 _1219_ (.A0(net96),
    .A1(\cpu_inst.IRHOLD[6] ),
    .S(net75),
    .X(_0648_));
 sky130_fd_sc_hd__nand2_2 _1220_ (.A(net49),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__inv_2 _1221_ (.A(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _1222_ (.A(_0620_),
    .B(_0649_),
    .Y(_0651_));
 sky130_fd_sc_hd__or2_1 _1223_ (.A(_0620_),
    .B(_0649_),
    .X(_0652_));
 sky130_fd_sc_hd__and2b_1 _1224_ (.A_N(net75),
    .B(\cpu_inst.DI[5] ),
    .X(_0653_));
 sky130_fd_sc_hd__a21oi_2 _1225_ (.A1(net75),
    .A2(\cpu_inst.IRHOLD[5] ),
    .B1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__a21o_2 _1226_ (.A1(\cpu_inst.IRHOLD_valid ),
    .A2(\cpu_inst.IRHOLD[5] ),
    .B1(_0653_),
    .X(_0655_));
 sky130_fd_sc_hd__and2_2 _1227_ (.A(net49),
    .B(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__nor3_1 _1228_ (.A(_0545_),
    .B(_0652_),
    .C(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__a31o_1 _1229_ (.A1(net30),
    .A2(_0646_),
    .A3(_0657_),
    .B1(_0642_),
    .X(_0658_));
 sky130_fd_sc_hd__o211a_1 _1230_ (.A1(net84),
    .A2(\cpu_inst.store ),
    .B1(net57),
    .C1(_0625_),
    .X(_0659_));
 sky130_fd_sc_hd__nor2_1 _1231_ (.A(_0562_),
    .B(_0639_),
    .Y(_0660_));
 sky130_fd_sc_hd__or4_1 _1232_ (.A(_0638_),
    .B(_0658_),
    .C(_0659_),
    .D(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__or2_1 _1233_ (.A(_0608_),
    .B(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(net54),
    .B(_0600_),
    .Y(_0663_));
 sky130_fd_sc_hd__nor2_2 _1235_ (.A(_0613_),
    .B(_0644_),
    .Y(_0664_));
 sky130_fd_sc_hd__or2_1 _1236_ (.A(_0613_),
    .B(_0644_),
    .X(_0665_));
 sky130_fd_sc_hd__or3_2 _1237_ (.A(_0545_),
    .B(_0656_),
    .C(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__nand2_1 _1238_ (.A(net29),
    .B(_0622_),
    .Y(_0667_));
 sky130_fd_sc_hd__nor2_1 _1239_ (.A(_0666_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__a21o_1 _1240_ (.A1(net68),
    .A2(_0663_),
    .B1(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__nor2_2 _1241_ (.A(net53),
    .B(_0639_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _1242_ (.A(net28),
    .B(_0546_),
    .Y(_0671_));
 sky130_fd_sc_hd__a22o_1 _1243_ (.A1(net70),
    .A2(net37),
    .B1(_0671_),
    .B2(_0646_),
    .X(_0672_));
 sky130_fd_sc_hd__nand2_2 _1244_ (.A(net86),
    .B(net85),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_1 _1245_ (.A(_0600_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__or4_4 _1246_ (.A(net94),
    .B(net91),
    .C(net87),
    .D(net89),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _1247_ (.A(_0673_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__mux2_1 _1248_ (.A0(_0674_),
    .A1(_0676_),
    .S(net58),
    .X(_0677_));
 sky130_fd_sc_hd__nor2_1 _1249_ (.A(\cpu_inst.state[5] ),
    .B(_0600_),
    .Y(_0678_));
 sky130_fd_sc_hd__and4bb_1 _1250_ (.A_N(net92),
    .B_N(net90),
    .C(net87),
    .D(net94),
    .X(_0679_));
 sky130_fd_sc_hd__or3b_2 _1251_ (.A(net90),
    .B(_0599_),
    .C_N(net87),
    .X(_0680_));
 sky130_fd_sc_hd__nor2_1 _1252_ (.A(net58),
    .B(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__or4b_4 _1253_ (.A(net93),
    .B(net91),
    .C(net89),
    .D_N(net88),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_1 _1254_ (.A(net70),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_1 _1255_ (.A(net86),
    .B(_0682_),
    .Y(_0684_));
 sky130_fd_sc_hd__or2_2 _1256_ (.A(\cpu_inst.state[4] ),
    .B(_0682_),
    .X(_0685_));
 sky130_fd_sc_hd__nor2_1 _1257_ (.A(net52),
    .B(_0682_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_2 _1258_ (.A(_0535_),
    .B(_0679_),
    .Y(_0687_));
 sky130_fd_sc_hd__o21a_1 _1259_ (.A1(_0681_),
    .A2(_0683_),
    .B1(_0673_),
    .X(_0688_));
 sky130_fd_sc_hd__nor2_1 _1260_ (.A(net85),
    .B(_0675_),
    .Y(_0689_));
 sky130_fd_sc_hd__mux2_1 _1261_ (.A0(_0678_),
    .A1(_0689_),
    .S(net58),
    .X(_0690_));
 sky130_fd_sc_hd__or2_1 _1262_ (.A(_0677_),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__or4_1 _1263_ (.A(_0669_),
    .B(_0672_),
    .C(_0688_),
    .D(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__or2_1 _1264_ (.A(_0662_),
    .B(_0692_),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _1265_ (.A(_0617_),
    .B(_0645_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _1266_ (.A0(_0604_),
    .A1(net38),
    .S(net68),
    .X(_0694_));
 sky130_fd_sc_hd__a21oi_1 _1267_ (.A1(net68),
    .A2(_0550_),
    .B1(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__o31a_1 _1268_ (.A1(net28),
    .A2(_0545_),
    .A3(_0693_),
    .B1(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_2 _1269_ (.A(_0544_),
    .B(_0656_),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_1 _1270_ (.A(_0644_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__nand2_1 _1271_ (.A(net68),
    .B(_0579_),
    .Y(_0699_));
 sky130_fd_sc_hd__o31a_1 _1272_ (.A1(_0665_),
    .A2(_0667_),
    .A3(_0697_),
    .B1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nand2_1 _1273_ (.A(_0696_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(net58),
    .B(_0568_),
    .Y(_0702_));
 sky130_fd_sc_hd__o221a_1 _1275_ (.A1(_0556_),
    .A2(_0562_),
    .B1(_0680_),
    .B2(_0561_),
    .C1(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__or3b_2 _1276_ (.A(_0611_),
    .B(_0644_),
    .C_N(_0531_),
    .X(_0704_));
 sky130_fd_sc_hd__nand2_1 _1277_ (.A(net30),
    .B(_0657_),
    .Y(_0705_));
 sky130_fd_sc_hd__o21ai_1 _1278_ (.A1(_0704_),
    .A2(_0705_),
    .B1(_0703_),
    .Y(_0706_));
 sky130_fd_sc_hd__mux4_2 _1279_ (.A0(\cpu_inst.N ),
    .A1(\cpu_inst.V ),
    .A2(\cpu_inst.C ),
    .A3(\cpu_inst.Z ),
    .S0(\cpu_inst.cond_code[1] ),
    .S1(\cpu_inst.cond_code[2] ),
    .X(_0707_));
 sky130_fd_sc_hd__xnor2_1 _1280_ (.A(\cpu_inst.cond_code[0] ),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__mux2_1 _1281_ (.A0(_0558_),
    .A1(_0640_),
    .S(net59),
    .X(_0709_));
 sky130_fd_sc_hd__a31o_1 _1282_ (.A1(net56),
    .A2(net37),
    .A3(_0708_),
    .B1(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__a2111o_1 _1283_ (.A1(net70),
    .A2(net42),
    .B1(_0701_),
    .C1(_0706_),
    .D1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__or2_1 _1284_ (.A(_0652_),
    .B(_0697_),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_1 _1285_ (.A(_0622_),
    .B(_0649_),
    .Y(_0713_));
 sky130_fd_sc_hd__inv_2 _1286_ (.A(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__or2_2 _1287_ (.A(_0697_),
    .B(_0713_),
    .X(_0715_));
 sky130_fd_sc_hd__o22a_1 _1288_ (.A1(_0562_),
    .A2(_0565_),
    .B1(_0647_),
    .B2(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__o221ai_2 _1289_ (.A1(net56),
    .A2(_0575_),
    .B1(_0647_),
    .B2(_0712_),
    .C1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__o32a_1 _1290_ (.A1(_0647_),
    .A2(_0652_),
    .A3(_0697_),
    .B1(_0575_),
    .B2(net56),
    .X(_0718_));
 sky130_fd_sc_hd__inv_2 _1291_ (.A(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__or2_1 _1292_ (.A(_0711_),
    .B(_0717_),
    .X(_0720_));
 sky130_fd_sc_hd__o32a_1 _1293_ (.A1(net28),
    .A2(_0546_),
    .A3(_0693_),
    .B1(_0586_),
    .B2(_0562_),
    .X(_0721_));
 sky130_fd_sc_hd__nor2_2 _1294_ (.A(net54),
    .B(_0586_),
    .Y(_0722_));
 sky130_fd_sc_hd__mux2_1 _1295_ (.A0(_0663_),
    .A1(_0722_),
    .S(net71),
    .X(_0723_));
 sky130_fd_sc_hd__nand2_1 _1296_ (.A(net59),
    .B(_0687_),
    .Y(_0724_));
 sky130_fd_sc_hd__o21a_1 _1297_ (.A1(net56),
    .A2(net46),
    .B1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__a21o_1 _1298_ (.A1(_0588_),
    .A2(_0724_),
    .B1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__o211a_1 _1299_ (.A1(_0531_),
    .A2(_0618_),
    .B1(_0671_),
    .C1(_0612_),
    .X(_0727_));
 sky130_fd_sc_hd__or4b_1 _1300_ (.A(_0723_),
    .B(_0726_),
    .C(_0727_),
    .D_N(_0721_),
    .X(_0728_));
 sky130_fd_sc_hd__or3_1 _1301_ (.A(_0608_),
    .B(_0720_),
    .C(_0728_),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _1302_ (.A(net55),
    .B(_0595_),
    .Y(_0729_));
 sky130_fd_sc_hd__or2_2 _1303_ (.A(net55),
    .B(_0595_),
    .X(_0730_));
 sky130_fd_sc_hd__nor2_2 _1304_ (.A(_0614_),
    .B(_0643_),
    .Y(_0731_));
 sky130_fd_sc_hd__or2_1 _1305_ (.A(_0614_),
    .B(_0643_),
    .X(_0732_));
 sky130_fd_sc_hd__o221a_1 _1306_ (.A1(_0544_),
    .A2(_0614_),
    .B1(_0622_),
    .B2(_0644_),
    .C1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__o32ai_4 _1307_ (.A1(net28),
    .A2(_0613_),
    .A3(_0733_),
    .B1(_0730_),
    .B2(net56),
    .Y(_0734_));
 sky130_fd_sc_hd__o311a_1 _1308_ (.A1(net84),
    .A2(\cpu_inst.write_back ),
    .A3(\cpu_inst.store ),
    .B1(net56),
    .C1(_0593_),
    .X(_0735_));
 sky130_fd_sc_hd__a211o_1 _1309_ (.A1(net68),
    .A2(_0596_),
    .B1(_0734_),
    .C1(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__or4_1 _1310_ (.A(_0564_),
    .B(_0585_),
    .C(_0672_),
    .D(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__or3_1 _1311_ (.A(net52),
    .B(_0556_),
    .C(_0583_),
    .X(_0738_));
 sky130_fd_sc_hd__o211a_1 _1312_ (.A1(net85),
    .A2(_0553_),
    .B1(_0635_),
    .C1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__a41o_1 _1313_ (.A1(_0586_),
    .A2(_0595_),
    .A3(_0675_),
    .A4(_0680_),
    .B1(net54),
    .X(_0740_));
 sky130_fd_sc_hd__a21o_1 _1314_ (.A1(_0739_),
    .A2(_0740_),
    .B1(net69),
    .X(_0741_));
 sky130_fd_sc_hd__or3b_1 _1315_ (.A(net70),
    .B(_0708_),
    .C_N(net37),
    .X(_0742_));
 sky130_fd_sc_hd__or2_1 _1316_ (.A(net54),
    .B(_0537_),
    .X(_0743_));
 sky130_fd_sc_hd__or2_1 _1317_ (.A(net69),
    .B(_0574_),
    .X(_0744_));
 sky130_fd_sc_hd__o21ai_1 _1318_ (.A1(net58),
    .A2(_0743_),
    .B1(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__or2_1 _1319_ (.A(_0537_),
    .B(net50),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _1320_ (.A0(_0572_),
    .A1(_0746_),
    .S(net69),
    .X(_0747_));
 sky130_fd_sc_hd__o311a_1 _1321_ (.A1(net86),
    .A2(net58),
    .A3(_0537_),
    .B1(_0744_),
    .C1(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__and3_1 _1322_ (.A(_0741_),
    .B(_0742_),
    .C(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__o22a_1 _1323_ (.A1(_0561_),
    .A2(_0589_),
    .B1(_0595_),
    .B2(_0562_),
    .X(_0750_));
 sky130_fd_sc_hd__nand2_1 _1324_ (.A(_0749_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__or4_1 _1325_ (.A(_0661_),
    .B(_0711_),
    .C(_0737_),
    .D(_0751_),
    .X(_0011_));
 sky130_fd_sc_hd__a22o_1 _1326_ (.A1(_0534_),
    .A2(_0671_),
    .B1(_0676_),
    .B2(net70),
    .X(_0752_));
 sky130_fd_sc_hd__a2bb2o_1 _1327_ (.A1_N(_0562_),
    .A2_N(_0675_),
    .B1(net56),
    .B2(_0548_),
    .X(_0753_));
 sky130_fd_sc_hd__nor2_1 _1328_ (.A(_0752_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__or2_2 _1329_ (.A(net71),
    .B(_0580_),
    .X(_0755_));
 sky130_fd_sc_hd__o21ai_1 _1330_ (.A1(net54),
    .A2(_0675_),
    .B1(net68),
    .Y(_0756_));
 sky130_fd_sc_hd__o21ai_1 _1331_ (.A1(net86),
    .A2(_0675_),
    .B1(net70),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2_1 _1332_ (.A(net59),
    .B(_0554_),
    .Y(_0758_));
 sky130_fd_sc_hd__o31a_1 _1333_ (.A1(_0500_),
    .A2(net56),
    .A3(_0685_),
    .B1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__o32a_1 _1334_ (.A1(net28),
    .A2(_0704_),
    .A3(_0712_),
    .B1(_0562_),
    .B2(_0682_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_1 _1335_ (.A(_0759_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__or2_1 _1336_ (.A(_0543_),
    .B(_0704_),
    .X(_0762_));
 sky130_fd_sc_hd__o2111ai_1 _1337_ (.A1(_0618_),
    .A2(_0731_),
    .B1(_0531_),
    .C1(_0544_),
    .D1(_0612_),
    .Y(_0763_));
 sky130_fd_sc_hd__o221a_1 _1338_ (.A1(_0704_),
    .A2(_0715_),
    .B1(_0762_),
    .B2(_0622_),
    .C1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__o21ai_1 _1339_ (.A1(net28),
    .A2(_0764_),
    .B1(_0754_),
    .Y(_0765_));
 sky130_fd_sc_hd__a2111o_1 _1340_ (.A1(_0755_),
    .A2(_0757_),
    .B1(_0765_),
    .C1(_0736_),
    .D1(_0692_),
    .X(_0766_));
 sky130_fd_sc_hd__or4_1 _1341_ (.A(_0728_),
    .B(_0751_),
    .C(_0761_),
    .D(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__or3_1 _1342_ (.A(_0662_),
    .B(_0720_),
    .C(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__or3_1 _1343_ (.A(_0577_),
    .B(_0581_),
    .C(_0725_),
    .X(_0769_));
 sky130_fd_sc_hd__or4b_1 _1344_ (.A(_0552_),
    .B(_0769_),
    .C(_0688_),
    .D_N(_0749_),
    .X(_0770_));
 sky130_fd_sc_hd__or4_1 _1345_ (.A(_0638_),
    .B(_0717_),
    .C(_0761_),
    .D(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__or3b_1 _1346_ (.A(_0701_),
    .B(_0771_),
    .C_N(_0768_),
    .X(_0012_));
 sky130_fd_sc_hd__a31o_1 _1347_ (.A1(net86),
    .A2(net67),
    .A3(_0689_),
    .B1(_0563_),
    .X(_0772_));
 sky130_fd_sc_hd__or4_1 _1348_ (.A(_0573_),
    .B(_0581_),
    .C(_0592_),
    .D(_0659_),
    .X(_0773_));
 sky130_fd_sc_hd__o311a_1 _1349_ (.A1(_0610_),
    .A2(_0681_),
    .A3(_0683_),
    .B1(_0500_),
    .C1(net86),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _1350_ (.A(_0747_),
    .B(_0750_),
    .Y(_0775_));
 sky130_fd_sc_hd__a2111o_1 _1351_ (.A1(net70),
    .A2(_0631_),
    .B1(_0677_),
    .C1(_0774_),
    .D1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__or3_1 _1352_ (.A(_0772_),
    .B(_0773_),
    .C(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _1353_ (.A(_0716_),
    .B(_0754_),
    .Y(_0778_));
 sky130_fd_sc_hd__and2_1 _1354_ (.A(_0700_),
    .B(_0760_),
    .X(_0779_));
 sky130_fd_sc_hd__and3b_1 _1355_ (.A_N(_0706_),
    .B(_0721_),
    .C(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__or3b_1 _1356_ (.A(_0777_),
    .B(_0778_),
    .C_N(_0780_),
    .X(_0013_));
 sky130_fd_sc_hd__o31a_1 _1357_ (.A1(_0610_),
    .A2(_0681_),
    .A3(_0683_),
    .B1(_0524_),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _1358_ (.A(_0559_),
    .B(_0576_),
    .Y(_0782_));
 sky130_fd_sc_hd__or4b_1 _1359_ (.A(_0606_),
    .B(_0719_),
    .C(_0781_),
    .D_N(_0759_),
    .X(_0783_));
 sky130_fd_sc_hd__a2111o_1 _1360_ (.A1(_0755_),
    .A2(_0756_),
    .B1(_0694_),
    .C1(_0709_),
    .D1(_0745_),
    .X(_0784_));
 sky130_fd_sc_hd__or4_1 _1361_ (.A(_0677_),
    .B(_0723_),
    .C(_0782_),
    .D(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__or4_1 _1362_ (.A(_0547_),
    .B(_0669_),
    .C(_0752_),
    .D(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__or4_1 _1363_ (.A(_0658_),
    .B(_0734_),
    .C(_0783_),
    .D(_0786_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _1364_ (.A(net209),
    .B(net226),
    .X(_0000_));
 sky130_fd_sc_hd__o21a_1 _1365_ (.A1(\spi_sram_master_inst.state[5] ),
    .A2(\spi_sram_master_inst.state[3] ),
    .B1(net207),
    .X(_0003_));
 sky130_fd_sc_hd__o21a_1 _1366_ (.A1(\spi_sram_master_inst.state[5] ),
    .A2(net221),
    .B1(_0506_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1367_ (.A(net223),
    .B(net226),
    .X(_0001_));
 sky130_fd_sc_hd__nand3_1 _1368_ (.A(net127),
    .B(_0511_),
    .C(_0518_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(net127),
    .B(net201),
    .Y(_0787_));
 sky130_fd_sc_hd__a21oi_1 _1370_ (.A1(_0512_),
    .A2(_0787_),
    .B1(_0521_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_2 _1371_ (.A(_0572_),
    .B(_0687_),
    .Y(_0788_));
 sky130_fd_sc_hd__nor2_1 _1372_ (.A(_0686_),
    .B(_0722_),
    .Y(_0789_));
 sky130_fd_sc_hd__o2111ai_4 _1373_ (.A1(\cpu_inst.state[5] ),
    .A2(_0565_),
    .B1(_0572_),
    .C1(_0687_),
    .D1(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_2 _1374_ (.A(_0632_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__or2_1 _1375_ (.A(net38),
    .B(_0790_),
    .X(_0792_));
 sky130_fd_sc_hd__nand3_1 _1376_ (.A(_0569_),
    .B(_0743_),
    .C(_0746_),
    .Y(_0793_));
 sky130_fd_sc_hd__nand2_1 _1377_ (.A(net44),
    .B(_0575_),
    .Y(_0794_));
 sky130_fd_sc_hd__or4_1 _1378_ (.A(_0579_),
    .B(_0580_),
    .C(_0684_),
    .D(_0722_),
    .X(_0795_));
 sky130_fd_sc_hd__nor4_1 _1379_ (.A(_0640_),
    .B(_0793_),
    .C(_0794_),
    .D(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__or4_2 _1380_ (.A(_0640_),
    .B(_0793_),
    .C(_0794_),
    .D(_0795_),
    .X(_0797_));
 sky130_fd_sc_hd__o22a_1 _1381_ (.A1(net53),
    .A2(_0549_),
    .B1(net51),
    .B2(_0589_),
    .X(_0798_));
 sky130_fd_sc_hd__o22a_1 _1382_ (.A1(net52),
    .A2(_0586_),
    .B1(_0673_),
    .B2(_0675_),
    .X(_0799_));
 sky130_fd_sc_hd__nand2_2 _1383_ (.A(_0798_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__and4_1 _1384_ (.A(\cpu_inst.src_reg[0] ),
    .B(net47),
    .C(_0798_),
    .D(_0799_),
    .X(_0801_));
 sky130_fd_sc_hd__a221o_1 _1385_ (.A1(\cpu_inst.dst_reg[0] ),
    .A2(net48),
    .B1(_0800_),
    .B2(\cpu_inst.index_y ),
    .C1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__nor2_1 _1386_ (.A(_0797_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__and2_1 _1387_ (.A(\cpu_inst.dst_reg[1] ),
    .B(net48),
    .X(_0804_));
 sky130_fd_sc_hd__a311oi_4 _1388_ (.A1(\cpu_inst.src_reg[1] ),
    .A2(net47),
    .A3(net20),
    .B1(_0800_),
    .C1(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__a311o_4 _1389_ (.A1(\cpu_inst.src_reg[1] ),
    .A2(net47),
    .A3(_0796_),
    .B1(_0800_),
    .C1(_0804_),
    .X(_0806_));
 sky130_fd_sc_hd__or3_1 _1390_ (.A(_0502_),
    .B(_0797_),
    .C(_0802_),
    .X(_0807_));
 sky130_fd_sc_hd__o211ai_1 _1391_ (.A1(_0503_),
    .A2(net16),
    .B1(_0806_),
    .C1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__or2_2 _1392_ (.A(net16),
    .B(_0806_),
    .X(_0809_));
 sky130_fd_sc_hd__o21a_1 _1393_ (.A1(_0797_),
    .A2(_0802_),
    .B1(\cpu_inst.AXYS[1][0] ),
    .X(_0810_));
 sky130_fd_sc_hd__a211o_1 _1394_ (.A1(\cpu_inst.AXYS[0][0] ),
    .A2(net16),
    .B1(_0806_),
    .C1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__and2_1 _1395_ (.A(_0808_),
    .B(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__o21ai_4 _1396_ (.A1(\cpu_inst.state[5] ),
    .A2(_0685_),
    .B1(net44),
    .Y(_0813_));
 sky130_fd_sc_hd__a21o_2 _1397_ (.A1(\cpu_inst.php ),
    .A2(_0722_),
    .B1(net45),
    .X(_0814_));
 sky130_fd_sc_hd__a21o_1 _1398_ (.A1(_0508_),
    .A2(_0722_),
    .B1(net38),
    .X(_0815_));
 sky130_fd_sc_hd__a22o_1 _1399_ (.A1(\cpu_inst.PC[0] ),
    .A2(_0788_),
    .B1(_0814_),
    .B2(\cpu_inst.C ),
    .X(_0816_));
 sky130_fd_sc_hd__a221o_1 _1400_ (.A1(\cpu_inst.PC[8] ),
    .A2(_0813_),
    .B1(_0815_),
    .B2(net83),
    .C1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__a211o_1 _1401_ (.A1(_0791_),
    .A2(_0812_),
    .B1(_0817_),
    .C1(net72),
    .X(_0818_));
 sky130_fd_sc_hd__or4_4 _1402_ (.A(\spi_sram_master_inst.state[1] ),
    .B(\spi_sram_master_inst.state[2] ),
    .C(\spi_sram_master_inst.state[6] ),
    .D(\spi_sram_master_inst.state[4] ),
    .X(_0819_));
 sky130_fd_sc_hd__nor2_1 _1403_ (.A(net61),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__or2_4 _1404_ (.A(net61),
    .B(_0819_),
    .X(_0821_));
 sky130_fd_sc_hd__nor2_2 _1405_ (.A(net60),
    .B(net32),
    .Y(_0822_));
 sky130_fd_sc_hd__nand2_2 _1406_ (.A(net71),
    .B(_0819_),
    .Y(_0823_));
 sky130_fd_sc_hd__o221a_1 _1407_ (.A1(net100),
    .A2(_0821_),
    .B1(_0823_),
    .B2(net4),
    .C1(_0818_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1408_ (.A0(\cpu_inst.AXYS[3][1] ),
    .A1(\cpu_inst.AXYS[2][1] ),
    .S(net17),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _1409_ (.A0(\cpu_inst.AXYS[1][1] ),
    .A1(\cpu_inst.AXYS[0][1] ),
    .S(net17),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_2 _1410_ (.A0(_0824_),
    .A1(_0825_),
    .S(net15),
    .X(_0826_));
 sky130_fd_sc_hd__or2_1 _1411_ (.A(net72),
    .B(_0814_),
    .X(_0827_));
 sky130_fd_sc_hd__a22o_1 _1412_ (.A1(\cpu_inst.PC[9] ),
    .A2(_0813_),
    .B1(_0815_),
    .B2(net82),
    .X(_0828_));
 sky130_fd_sc_hd__a221o_1 _1413_ (.A1(\cpu_inst.PC[1] ),
    .A2(_0788_),
    .B1(_0814_),
    .B2(\cpu_inst.Z ),
    .C1(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__a211o_1 _1414_ (.A1(_0791_),
    .A2(_0826_),
    .B1(_0829_),
    .C1(net72),
    .X(_0830_));
 sky130_fd_sc_hd__a21o_1 _1415_ (.A1(net100),
    .A2(_0819_),
    .B1(net62),
    .X(_0831_));
 sky130_fd_sc_hd__a22o_1 _1416_ (.A1(net175),
    .A2(net35),
    .B1(_0830_),
    .B2(_0831_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1417_ (.A0(\cpu_inst.AXYS[3][2] ),
    .A1(\cpu_inst.AXYS[2][2] ),
    .S(net17),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _1418_ (.A0(\cpu_inst.AXYS[1][2] ),
    .A1(\cpu_inst.AXYS[0][2] ),
    .S(net17),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_2 _1419_ (.A0(_0832_),
    .A1(_0833_),
    .S(net15),
    .X(_0834_));
 sky130_fd_sc_hd__a22o_1 _1420_ (.A1(\cpu_inst.PC[10] ),
    .A2(_0813_),
    .B1(_0815_),
    .B2(net81),
    .X(_0835_));
 sky130_fd_sc_hd__a221o_1 _1421_ (.A1(\cpu_inst.PC[2] ),
    .A2(_0788_),
    .B1(_0814_),
    .B2(\cpu_inst.I ),
    .C1(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__a211o_1 _1422_ (.A1(_0791_),
    .A2(_0834_),
    .B1(_0836_),
    .C1(net72),
    .X(_0837_));
 sky130_fd_sc_hd__a21o_1 _1423_ (.A1(net99),
    .A2(_0819_),
    .B1(net62),
    .X(_0838_));
 sky130_fd_sc_hd__a22o_1 _1424_ (.A1(net98),
    .A2(net35),
    .B1(_0837_),
    .B2(_0838_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1425_ (.A0(\cpu_inst.AXYS[1][3] ),
    .A1(\cpu_inst.AXYS[0][3] ),
    .S(net17),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _1426_ (.A0(\cpu_inst.AXYS[3][3] ),
    .A1(\cpu_inst.AXYS[2][3] ),
    .S(net17),
    .X(_0840_));
 sky130_fd_sc_hd__or2_1 _1427_ (.A(net15),
    .B(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__o21ai_2 _1428_ (.A1(_0806_),
    .A2(_0839_),
    .B1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__nor2_1 _1429_ (.A(_0792_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__a221o_1 _1430_ (.A1(\cpu_inst.PC[3] ),
    .A2(_0788_),
    .B1(_0813_),
    .B2(\cpu_inst.PC[11] ),
    .C1(net72),
    .X(_0844_));
 sky130_fd_sc_hd__a221o_1 _1431_ (.A1(\cpu_inst.D ),
    .A2(_0814_),
    .B1(_0815_),
    .B2(net80),
    .C1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__o22a_1 _1432_ (.A1(net98),
    .A2(net63),
    .B1(_0843_),
    .B2(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _1433_ (.A0(net97),
    .A1(_0846_),
    .S(_0821_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(\cpu_inst.AXYS[1][4] ),
    .A1(\cpu_inst.AXYS[0][4] ),
    .S(net17),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _1435_ (.A0(\cpu_inst.AXYS[3][4] ),
    .A1(\cpu_inst.AXYS[2][4] ),
    .S(net17),
    .X(_0848_));
 sky130_fd_sc_hd__or2_1 _1436_ (.A(net15),
    .B(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__o21ai_2 _1437_ (.A1(_0806_),
    .A2(_0847_),
    .B1(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__nor2_1 _1438_ (.A(_0792_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__o21a_1 _1439_ (.A1(net38),
    .A2(_0722_),
    .B1(net79),
    .X(_0852_));
 sky130_fd_sc_hd__a221o_1 _1440_ (.A1(\cpu_inst.php ),
    .A2(_0722_),
    .B1(_0788_),
    .B2(\cpu_inst.PC[4] ),
    .C1(net72),
    .X(_0853_));
 sky130_fd_sc_hd__a221o_1 _1441_ (.A1(_0529_),
    .A2(net45),
    .B1(_0813_),
    .B2(\cpu_inst.PC[12] ),
    .C1(_0852_),
    .X(_0854_));
 sky130_fd_sc_hd__or3_1 _1442_ (.A(_0851_),
    .B(_0853_),
    .C(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__o221a_1 _1443_ (.A1(\cpu_inst.DI[4] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(net97),
    .C1(_0855_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(\cpu_inst.AXYS[1][5] ),
    .A1(\cpu_inst.AXYS[0][5] ),
    .S(net16),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(\cpu_inst.AXYS[3][5] ),
    .A1(\cpu_inst.AXYS[2][5] ),
    .S(net16),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_2 _1446_ (.A0(_0856_),
    .A1(_0857_),
    .S(_0806_),
    .X(_0858_));
 sky130_fd_sc_hd__o21a_1 _1447_ (.A1(net38),
    .A2(_0722_),
    .B1(net78),
    .X(_0859_));
 sky130_fd_sc_hd__a221o_1 _1448_ (.A1(\cpu_inst.PC[5] ),
    .A2(_0788_),
    .B1(_0813_),
    .B2(\cpu_inst.PC[13] ),
    .C1(_0827_),
    .X(_0860_));
 sky130_fd_sc_hd__a211o_1 _1449_ (.A1(_0791_),
    .A2(_0858_),
    .B1(_0859_),
    .C1(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__o221a_1 _1450_ (.A1(\cpu_inst.DI[5] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(\cpu_inst.DI[4] ),
    .C1(_0861_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(\cpu_inst.AXYS[1][6] ),
    .A1(\cpu_inst.AXYS[0][6] ),
    .S(net17),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(\cpu_inst.AXYS[3][6] ),
    .A1(\cpu_inst.AXYS[2][6] ),
    .S(net17),
    .X(_0863_));
 sky130_fd_sc_hd__or2_1 _1453_ (.A(net15),
    .B(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__o21ai_2 _1454_ (.A1(_0806_),
    .A2(_0862_),
    .B1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__nor2_1 _1455_ (.A(_0792_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__a221o_1 _1456_ (.A1(\cpu_inst.PC[6] ),
    .A2(_0788_),
    .B1(_0813_),
    .B2(\cpu_inst.PC[14] ),
    .C1(net72),
    .X(_0867_));
 sky130_fd_sc_hd__a22o_1 _1457_ (.A1(\cpu_inst.V ),
    .A2(_0814_),
    .B1(_0815_),
    .B2(net77),
    .X(_0868_));
 sky130_fd_sc_hd__o32a_1 _1458_ (.A1(_0866_),
    .A2(_0867_),
    .A3(_0868_),
    .B1(net63),
    .B2(\cpu_inst.DI[5] ),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _1459_ (.A0(net96),
    .A1(_0869_),
    .S(_0821_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1460_ (.A0(\cpu_inst.AXYS[1][7] ),
    .A1(\cpu_inst.AXYS[0][7] ),
    .S(net16),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(\cpu_inst.AXYS[3][7] ),
    .A1(\cpu_inst.AXYS[2][7] ),
    .S(net16),
    .X(_0871_));
 sky130_fd_sc_hd__or2_1 _1462_ (.A(net15),
    .B(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__o21ai_2 _1463_ (.A1(_0806_),
    .A2(_0870_),
    .B1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_1 _1464_ (.A(_0792_),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__a221o_1 _1465_ (.A1(\cpu_inst.PC[7] ),
    .A2(_0788_),
    .B1(_0813_),
    .B2(\cpu_inst.PC[15] ),
    .C1(net72),
    .X(_0875_));
 sky130_fd_sc_hd__a221o_1 _1466_ (.A1(\cpu_inst.N ),
    .A2(_0814_),
    .B1(_0815_),
    .B2(net76),
    .C1(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__o22a_1 _1467_ (.A1(net96),
    .A2(net63),
    .B1(_0874_),
    .B2(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(net95),
    .A1(_0877_),
    .S(_0821_),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _1469_ (.A(_0641_),
    .B(_0789_),
    .Y(_0878_));
 sky130_fd_sc_hd__nor2_1 _1470_ (.A(_0794_),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__or2_4 _1471_ (.A(_0794_),
    .B(_0878_),
    .X(_0880_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(_0557_),
    .B(_0687_),
    .Y(_0881_));
 sky130_fd_sc_hd__nand2_1 _1473_ (.A(_0572_),
    .B(_0574_),
    .Y(_0882_));
 sky130_fd_sc_hd__or3_1 _1474_ (.A(net46),
    .B(_0881_),
    .C(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__or3_4 _1475_ (.A(_0548_),
    .B(_0554_),
    .C(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__a2bb2o_1 _1476_ (.A1_N(_0553_),
    .A2_N(net51),
    .B1(_0601_),
    .B2(_0679_),
    .X(_0885_));
 sky130_fd_sc_hd__or3_4 _1477_ (.A(_0627_),
    .B(_0678_),
    .C(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__a21oi_1 _1478_ (.A1(_0537_),
    .A2(_0682_),
    .B1(net54),
    .Y(_0887_));
 sky130_fd_sc_hd__or2_1 _1479_ (.A(_0580_),
    .B(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__a2111o_1 _1480_ (.A1(\cpu_inst.state[4] ),
    .A2(_0689_),
    .B1(_0888_),
    .C1(_0591_),
    .D1(_0674_),
    .X(_0889_));
 sky130_fd_sc_hd__or3_4 _1481_ (.A(_0884_),
    .B(_0886_),
    .C(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__a211o_4 _1482_ (.A1(net90),
    .A2(_0631_),
    .B1(_0596_),
    .C1(net43),
    .X(_0891_));
 sky130_fd_sc_hd__or2_1 _1483_ (.A(_0604_),
    .B(_0729_),
    .X(_0892_));
 sky130_fd_sc_hd__or2_4 _1484_ (.A(net38),
    .B(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__or2_4 _1485_ (.A(_0891_),
    .B(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__or2_4 _1486_ (.A(_0528_),
    .B(_0590_),
    .X(_0895_));
 sky130_fd_sc_hd__or2_1 _1487_ (.A(net39),
    .B(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__nor4_1 _1488_ (.A(_0880_),
    .B(_0890_),
    .C(_0894_),
    .D(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__or4_4 _1489_ (.A(_0880_),
    .B(_0890_),
    .C(_0894_),
    .D(_0896_),
    .X(_0898_));
 sky130_fd_sc_hd__and2_1 _1490_ (.A(net83),
    .B(net40),
    .X(_0899_));
 sky130_fd_sc_hd__a221o_1 _1491_ (.A1(\cpu_inst.ABL[0] ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(net100),
    .C1(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__a221o_1 _1492_ (.A1(_0812_),
    .A2(_0880_),
    .B1(_0890_),
    .B2(net83),
    .C1(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(\cpu_inst.PC[0] ),
    .A1(_0901_),
    .S(_0898_),
    .X(_0902_));
 sky130_fd_sc_hd__a22o_1 _1494_ (.A1(net255),
    .A2(net36),
    .B1(net25),
    .B2(net95),
    .X(_0903_));
 sky130_fd_sc_hd__a21o_1 _1495_ (.A1(net64),
    .A2(_0902_),
    .B1(_0903_),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_1 _1496_ (.A1(net82),
    .A2(net39),
    .B1(_0895_),
    .B2(net99),
    .X(_0904_));
 sky130_fd_sc_hd__a211o_1 _1497_ (.A1(\cpu_inst.ABL[1] ),
    .A2(_0894_),
    .B1(net7),
    .C1(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__a22o_1 _1498_ (.A1(_0826_),
    .A2(_0880_),
    .B1(_0890_),
    .B2(net82),
    .X(_0906_));
 sky130_fd_sc_hd__o22a_1 _1499_ (.A1(\cpu_inst.PC[1] ),
    .A2(_0898_),
    .B1(_0905_),
    .B2(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__a22o_1 _1500_ (.A1(\spi_sram_master_inst.data[9] ),
    .A2(net35),
    .B1(net25),
    .B2(net255),
    .X(_0908_));
 sky130_fd_sc_hd__a21o_1 _1501_ (.A1(net64),
    .A2(_0907_),
    .B1(net256),
    .X(_0028_));
 sky130_fd_sc_hd__a22o_1 _1502_ (.A1(net81),
    .A2(net39),
    .B1(_0895_),
    .B2(net98),
    .X(_0909_));
 sky130_fd_sc_hd__a211o_1 _1503_ (.A1(\cpu_inst.ABL[2] ),
    .A2(_0894_),
    .B1(net7),
    .C1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _1504_ (.A1(_0834_),
    .A2(_0880_),
    .B1(_0890_),
    .B2(net81),
    .X(_0911_));
 sky130_fd_sc_hd__o22a_1 _1505_ (.A1(\cpu_inst.PC[2] ),
    .A2(_0898_),
    .B1(_0910_),
    .B2(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__a22o_1 _1506_ (.A1(net280),
    .A2(net35),
    .B1(net25),
    .B2(net262),
    .X(_0913_));
 sky130_fd_sc_hd__a21o_1 _1507_ (.A1(net64),
    .A2(_0912_),
    .B1(_0913_),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _1508_ (.A1(net80),
    .A2(net39),
    .B1(_0895_),
    .B2(net97),
    .X(_0914_));
 sky130_fd_sc_hd__a211o_1 _1509_ (.A1(\cpu_inst.ABL[3] ),
    .A2(_0894_),
    .B1(net7),
    .C1(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a2bb2o_1 _1510_ (.A1_N(_0842_),
    .A2_N(_0879_),
    .B1(_0890_),
    .B2(net80),
    .X(_0916_));
 sky130_fd_sc_hd__o22a_1 _1511_ (.A1(\cpu_inst.PC[3] ),
    .A2(_0898_),
    .B1(_0915_),
    .B2(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__a22o_1 _1512_ (.A1(net283),
    .A2(net35),
    .B1(net25),
    .B2(net265),
    .X(_0918_));
 sky130_fd_sc_hd__a21o_1 _1513_ (.A1(net64),
    .A2(_0917_),
    .B1(_0918_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _1514_ (.A1(net79),
    .A2(net39),
    .B1(_0895_),
    .B2(\cpu_inst.DI[4] ),
    .X(_0919_));
 sky130_fd_sc_hd__a211o_1 _1515_ (.A1(\cpu_inst.ABL[4] ),
    .A2(_0894_),
    .B1(net8),
    .C1(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__a2bb2o_1 _1516_ (.A1_N(_0850_),
    .A2_N(_0879_),
    .B1(_0890_),
    .B2(net79),
    .X(_0921_));
 sky130_fd_sc_hd__o22a_1 _1517_ (.A1(\cpu_inst.PC[4] ),
    .A2(_0898_),
    .B1(_0920_),
    .B2(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__a22o_1 _1518_ (.A1(net251),
    .A2(net35),
    .B1(net25),
    .B2(net278),
    .X(_0923_));
 sky130_fd_sc_hd__a21o_1 _1519_ (.A1(net64),
    .A2(_0922_),
    .B1(_0923_),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _1520_ (.A1(net78),
    .A2(net39),
    .B1(_0895_),
    .B2(\cpu_inst.DI[5] ),
    .X(_0924_));
 sky130_fd_sc_hd__a211o_1 _1521_ (.A1(\cpu_inst.ABL[5] ),
    .A2(_0894_),
    .B1(net8),
    .C1(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__a22o_1 _1522_ (.A1(_0858_),
    .A2(_0880_),
    .B1(_0890_),
    .B2(net78),
    .X(_0926_));
 sky130_fd_sc_hd__o22a_1 _1523_ (.A1(\cpu_inst.PC[5] ),
    .A2(_0898_),
    .B1(_0925_),
    .B2(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__a22o_1 _1524_ (.A1(\spi_sram_master_inst.data[13] ),
    .A2(net36),
    .B1(net25),
    .B2(net251),
    .X(_0928_));
 sky130_fd_sc_hd__a21o_1 _1525_ (.A1(net64),
    .A2(_0927_),
    .B1(net252),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _1526_ (.A1(net77),
    .A2(net39),
    .B1(_0895_),
    .B2(net96),
    .X(_0929_));
 sky130_fd_sc_hd__a211o_1 _1527_ (.A1(\cpu_inst.ABL[6] ),
    .A2(_0894_),
    .B1(net8),
    .C1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__a2bb2o_1 _1528_ (.A1_N(_0865_),
    .A2_N(_0879_),
    .B1(_0890_),
    .B2(net77),
    .X(_0931_));
 sky130_fd_sc_hd__o22a_1 _1529_ (.A1(\cpu_inst.PC[6] ),
    .A2(_0898_),
    .B1(_0930_),
    .B2(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__a22o_1 _1530_ (.A1(\spi_sram_master_inst.data[14] ),
    .A2(net36),
    .B1(_0822_),
    .B2(net263),
    .X(_0933_));
 sky130_fd_sc_hd__a21o_1 _1531_ (.A1(net64),
    .A2(_0932_),
    .B1(net264),
    .X(_0033_));
 sky130_fd_sc_hd__nor2_1 _1532_ (.A(_0873_),
    .B(_0879_),
    .Y(_0934_));
 sky130_fd_sc_hd__a221o_1 _1533_ (.A1(net76),
    .A2(_0890_),
    .B1(_0895_),
    .B2(net95),
    .C1(net8),
    .X(_0935_));
 sky130_fd_sc_hd__a221o_1 _1534_ (.A1(\cpu_inst.ADD[7] ),
    .A2(net39),
    .B1(_0894_),
    .B2(\cpu_inst.ABL[7] ),
    .C1(_0934_),
    .X(_0936_));
 sky130_fd_sc_hd__o22a_1 _1535_ (.A1(\cpu_inst.PC[7] ),
    .A2(_0898_),
    .B1(_0935_),
    .B2(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__a22o_1 _1536_ (.A1(\spi_sram_master_inst.data[15] ),
    .A2(net36),
    .B1(_0822_),
    .B2(net268),
    .X(_0938_));
 sky130_fd_sc_hd__a21o_1 _1537_ (.A1(net62),
    .A2(_0937_),
    .B1(_0938_),
    .X(_0034_));
 sky130_fd_sc_hd__a221o_1 _1538_ (.A1(net83),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[0] ),
    .C1(_0883_),
    .X(_0939_));
 sky130_fd_sc_hd__and2_1 _1539_ (.A(\cpu_inst.ABH[0] ),
    .B(net41),
    .X(_0940_));
 sky130_fd_sc_hd__or4_1 _1540_ (.A(_0554_),
    .B(_0880_),
    .C(_0888_),
    .D(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__a211o_1 _1541_ (.A1(net100),
    .A2(_0886_),
    .B1(_0939_),
    .C1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__a21o_1 _1542_ (.A1(\cpu_inst.PC[8] ),
    .A2(net7),
    .B1(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__a22o_1 _1543_ (.A1(net275),
    .A2(net35),
    .B1(net25),
    .B2(\spi_sram_master_inst.data[15] ),
    .X(_0944_));
 sky130_fd_sc_hd__a21o_1 _1544_ (.A1(net66),
    .A2(_0943_),
    .B1(net276),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _1545_ (.A(\cpu_inst.ABH[1] ),
    .B(net41),
    .X(_0945_));
 sky130_fd_sc_hd__a221o_1 _1546_ (.A1(net82),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[1] ),
    .C1(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__a221o_1 _1547_ (.A1(net99),
    .A2(_0886_),
    .B1(net7),
    .B2(\cpu_inst.PC[9] ),
    .C1(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__a22o_1 _1548_ (.A1(\spi_sram_master_inst.data[17] ),
    .A2(net35),
    .B1(net25),
    .B2(net281),
    .X(_0948_));
 sky130_fd_sc_hd__a21o_1 _1549_ (.A1(net62),
    .A2(_0947_),
    .B1(net282),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _1550_ (.A(\cpu_inst.ABH[2] ),
    .B(net41),
    .X(_0949_));
 sky130_fd_sc_hd__a221o_1 _1551_ (.A1(net81),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[2] ),
    .C1(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__a221o_1 _1552_ (.A1(net98),
    .A2(_0886_),
    .B1(net8),
    .B2(\cpu_inst.PC[10] ),
    .C1(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__a22o_1 _1553_ (.A1(\spi_sram_master_inst.data[18] ),
    .A2(net35),
    .B1(net25),
    .B2(net249),
    .X(_0952_));
 sky130_fd_sc_hd__a21o_1 _1554_ (.A1(net62),
    .A2(_0951_),
    .B1(_0952_),
    .X(_0037_));
 sky130_fd_sc_hd__and2_1 _1555_ (.A(\cpu_inst.ABH[3] ),
    .B(net41),
    .X(_0953_));
 sky130_fd_sc_hd__a221o_1 _1556_ (.A1(net80),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[3] ),
    .C1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__a221o_1 _1557_ (.A1(net97),
    .A2(_0886_),
    .B1(net7),
    .B2(\cpu_inst.PC[11] ),
    .C1(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__a22o_1 _1558_ (.A1(net272),
    .A2(net35),
    .B1(net25),
    .B2(\spi_sram_master_inst.data[18] ),
    .X(_0956_));
 sky130_fd_sc_hd__a21o_1 _1559_ (.A1(net62),
    .A2(_0955_),
    .B1(net273),
    .X(_0038_));
 sky130_fd_sc_hd__and2_1 _1560_ (.A(\cpu_inst.ABH[4] ),
    .B(net41),
    .X(_0957_));
 sky130_fd_sc_hd__a221o_1 _1561_ (.A1(net79),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[4] ),
    .C1(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__a221o_1 _1562_ (.A1(\cpu_inst.DI[4] ),
    .A2(_0886_),
    .B1(net7),
    .B2(\cpu_inst.PC[12] ),
    .C1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _1563_ (.A1(net260),
    .A2(net34),
    .B1(net24),
    .B2(\spi_sram_master_inst.data[19] ),
    .X(_0960_));
 sky130_fd_sc_hd__a21o_1 _1564_ (.A1(net62),
    .A2(_0959_),
    .B1(net261),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _1565_ (.A(\cpu_inst.ABH[5] ),
    .B(net41),
    .X(_0961_));
 sky130_fd_sc_hd__a221o_1 _1566_ (.A1(net78),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[5] ),
    .C1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__a221o_1 _1567_ (.A1(\cpu_inst.DI[5] ),
    .A2(_0886_),
    .B1(net7),
    .B2(\cpu_inst.PC[13] ),
    .C1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__a22o_1 _1568_ (.A1(\spi_sram_master_inst.data[21] ),
    .A2(net34),
    .B1(net24),
    .B2(net258),
    .X(_0964_));
 sky130_fd_sc_hd__a21o_1 _1569_ (.A1(net60),
    .A2(_0963_),
    .B1(net259),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _1570_ (.A(\cpu_inst.ABH[6] ),
    .B(net42),
    .X(_0965_));
 sky130_fd_sc_hd__a221o_1 _1571_ (.A1(net77),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[6] ),
    .C1(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__a221o_1 _1572_ (.A1(net96),
    .A2(_0886_),
    .B1(net7),
    .B2(\cpu_inst.PC[14] ),
    .C1(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__a22o_1 _1573_ (.A1(\spi_sram_master_inst.data[22] ),
    .A2(net34),
    .B1(net24),
    .B2(net266),
    .X(_0968_));
 sky130_fd_sc_hd__a21o_1 _1574_ (.A1(net60),
    .A2(_0967_),
    .B1(net267),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _1575_ (.A(\cpu_inst.ABH[7] ),
    .B(net42),
    .X(_0969_));
 sky130_fd_sc_hd__a221o_1 _1576_ (.A1(net76),
    .A2(_0891_),
    .B1(_0893_),
    .B2(\cpu_inst.ABH[7] ),
    .C1(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__a221o_1 _1577_ (.A1(net95),
    .A2(_0886_),
    .B1(net7),
    .B2(\cpu_inst.PC[15] ),
    .C1(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__a22o_1 _1578_ (.A1(net168),
    .A2(net34),
    .B1(net24),
    .B2(net271),
    .X(_0972_));
 sky130_fd_sc_hd__a21o_1 _1579_ (.A1(net60),
    .A2(_0971_),
    .B1(_0972_),
    .X(_0042_));
 sky130_fd_sc_hd__o21ai_1 _1580_ (.A1(_0603_),
    .A2(_0631_),
    .B1(\cpu_inst.store ),
    .Y(_0973_));
 sky130_fd_sc_hd__a21o_1 _1581_ (.A1(_0791_),
    .A2(_0973_),
    .B1(_0522_),
    .X(_0974_));
 sky130_fd_sc_hd__o221a_1 _1582_ (.A1(net165),
    .A2(_0821_),
    .B1(_0823_),
    .B2(net215),
    .C1(_0974_),
    .X(_0043_));
 sky130_fd_sc_hd__or3b_1 _1583_ (.A(net47),
    .B(net74),
    .C_N(\cpu_inst.load_reg ),
    .X(_0975_));
 sky130_fd_sc_hd__and3b_1 _1584_ (.A_N(_0888_),
    .B(_0746_),
    .C(_0569_),
    .X(_0976_));
 sky130_fd_sc_hd__a31o_2 _1585_ (.A1(net44),
    .A2(_0975_),
    .A3(_0976_),
    .B1(net71),
    .X(_0977_));
 sky130_fd_sc_hd__inv_2 _1586_ (.A(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__or3b_4 _1587_ (.A(_0805_),
    .B(_0977_),
    .C_N(net16),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _1588_ (.A0(\cpu_inst.DI[0] ),
    .A1(net83),
    .S(net44),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _1589_ (.A0(_0980_),
    .A1(net219),
    .S(_0979_),
    .X(_0044_));
 sky130_fd_sc_hd__and3_1 _1590_ (.A(\cpu_inst.adc_bcd ),
    .B(\cpu_inst.adj_bcd ),
    .C(\cpu_inst.ALU.HC ),
    .X(_0981_));
 sky130_fd_sc_hd__nand2b_1 _1591_ (.A_N(\cpu_inst.adc_bcd ),
    .B(\cpu_inst.adj_bcd ),
    .Y(_0982_));
 sky130_fd_sc_hd__nor2_1 _1592_ (.A(\cpu_inst.ALU.HC ),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__o21a_1 _1593_ (.A1(_0981_),
    .A2(_0983_),
    .B1(net82),
    .X(_0984_));
 sky130_fd_sc_hd__nor3_1 _1594_ (.A(net82),
    .B(_0981_),
    .C(_0983_),
    .Y(_0985_));
 sky130_fd_sc_hd__nor2_1 _1595_ (.A(_0984_),
    .B(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__mux2_1 _1596_ (.A0(net99),
    .A1(_0986_),
    .S(net44),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _1597_ (.A0(_0987_),
    .A1(net186),
    .S(_0979_),
    .X(_0045_));
 sky130_fd_sc_hd__nand2_1 _1598_ (.A(\cpu_inst.ADD[2] ),
    .B(_0981_),
    .Y(_0988_));
 sky130_fd_sc_hd__or2_1 _1599_ (.A(\cpu_inst.ADD[2] ),
    .B(_0981_),
    .X(_0989_));
 sky130_fd_sc_hd__nand2_1 _1600_ (.A(_0988_),
    .B(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__xnor2_1 _1601_ (.A(_0984_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__mux2_1 _1602_ (.A0(\cpu_inst.DI[2] ),
    .A1(_0991_),
    .S(net44),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _1603_ (.A0(_0992_),
    .A1(net185),
    .S(_0979_),
    .X(_0046_));
 sky130_fd_sc_hd__a21bo_1 _1604_ (.A1(_0984_),
    .A2(_0989_),
    .B1_N(_0988_),
    .X(_0993_));
 sky130_fd_sc_hd__xnor2_1 _1605_ (.A(\cpu_inst.ADD[3] ),
    .B(_0983_),
    .Y(_0994_));
 sky130_fd_sc_hd__xnor2_1 _1606_ (.A(_0993_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(\cpu_inst.DI[3] ),
    .A1(_0995_),
    .S(net44),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(_0996_),
    .A1(net172),
    .S(_0979_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(\cpu_inst.DI[4] ),
    .A1(\cpu_inst.ADD[4] ),
    .S(net44),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(_0997_),
    .A1(net193),
    .S(_0979_),
    .X(_0048_));
 sky130_fd_sc_hd__and3_1 _1611_ (.A(net84),
    .B(\cpu_inst.adc_bcd ),
    .C(\cpu_inst.adj_bcd ),
    .X(_0998_));
 sky130_fd_sc_hd__nor2_1 _1612_ (.A(net84),
    .B(_0982_),
    .Y(_0999_));
 sky130_fd_sc_hd__o21a_1 _1613_ (.A1(_0998_),
    .A2(_0999_),
    .B1(net78),
    .X(_1000_));
 sky130_fd_sc_hd__nor3_1 _1614_ (.A(net78),
    .B(_0998_),
    .C(_0999_),
    .Y(_1001_));
 sky130_fd_sc_hd__nor2_1 _1615_ (.A(_1000_),
    .B(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(\cpu_inst.DI[5] ),
    .A1(_1002_),
    .S(net44),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _1617_ (.A0(_1003_),
    .A1(net181),
    .S(_0979_),
    .X(_0049_));
 sky130_fd_sc_hd__nand2_1 _1618_ (.A(\cpu_inst.ADD[6] ),
    .B(_0998_),
    .Y(_1004_));
 sky130_fd_sc_hd__or2_1 _1619_ (.A(\cpu_inst.ADD[6] ),
    .B(_0998_),
    .X(_1005_));
 sky130_fd_sc_hd__nand2_1 _1620_ (.A(_1004_),
    .B(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__xnor2_1 _1621_ (.A(_1000_),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(\cpu_inst.DI[6] ),
    .A1(_1007_),
    .S(net44),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(_1008_),
    .A1(net189),
    .S(_0979_),
    .X(_0050_));
 sky130_fd_sc_hd__a21bo_1 _1624_ (.A1(_1000_),
    .A2(_1005_),
    .B1_N(_1004_),
    .X(_1009_));
 sky130_fd_sc_hd__xnor2_1 _1625_ (.A(\cpu_inst.ADD[7] ),
    .B(_0999_),
    .Y(_1010_));
 sky130_fd_sc_hd__xnor2_1 _1626_ (.A(_1009_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__mux2_1 _1627_ (.A0(\cpu_inst.DI[7] ),
    .A1(_1011_),
    .S(_0571_),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _1628_ (.A0(_1012_),
    .A1(net180),
    .S(_0979_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1629_ (.A0(net95),
    .A1(\cpu_inst.backwards ),
    .S(net71),
    .X(_0052_));
 sky130_fd_sc_hd__or2_4 _1630_ (.A(_0634_),
    .B(_0892_),
    .X(_1013_));
 sky130_fd_sc_hd__a221o_1 _1631_ (.A1(\cpu_inst.backwards ),
    .A2(net41),
    .B1(_1013_),
    .B2(\cpu_inst.op[2] ),
    .C1(_0790_),
    .X(_1014_));
 sky130_fd_sc_hd__and2_2 _1632_ (.A(\cpu_inst.op[3] ),
    .B(_1013_),
    .X(_1015_));
 sky130_fd_sc_hd__nand2_2 _1633_ (.A(\cpu_inst.op[3] ),
    .B(_1013_),
    .Y(_1016_));
 sky130_fd_sc_hd__or2_4 _1634_ (.A(_0604_),
    .B(net37),
    .X(_1017_));
 sky130_fd_sc_hd__nor2_1 _1635_ (.A(net46),
    .B(net42),
    .Y(_1018_));
 sky130_fd_sc_hd__or4b_1 _1636_ (.A(_0794_),
    .B(_0881_),
    .C(_1017_),
    .D_N(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__and2_1 _1637_ (.A(_0730_),
    .B(_0746_),
    .X(_1020_));
 sky130_fd_sc_hd__or3b_1 _1638_ (.A(_0663_),
    .B(_0882_),
    .C_N(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__or3_1 _1639_ (.A(_0548_),
    .B(_0554_),
    .C(_0579_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _1640_ (.A(_0558_),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__nor4b_2 _1641_ (.A(_0878_),
    .B(_1019_),
    .C(_1021_),
    .D_N(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__a22o_1 _1642_ (.A1(\cpu_inst.PC[6] ),
    .A2(net37),
    .B1(_1024_),
    .B2(net96),
    .X(_1025_));
 sky130_fd_sc_hd__or2_1 _1643_ (.A(_1015_),
    .B(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__xnor2_1 _1644_ (.A(net14),
    .B(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__or2_2 _1645_ (.A(_0579_),
    .B(_0663_),
    .X(_1028_));
 sky130_fd_sc_hd__o21ai_1 _1646_ (.A1(\cpu_inst.load_only ),
    .A2(_0635_),
    .B1(_1020_),
    .Y(_1029_));
 sky130_fd_sc_hd__or4_4 _1647_ (.A(_0800_),
    .B(_0880_),
    .C(_1028_),
    .D(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__inv_2 _1648_ (.A(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__a221o_1 _1649_ (.A1(net77),
    .A2(_0884_),
    .B1(_1017_),
    .B2(net96),
    .C1(_0965_),
    .X(_1032_));
 sky130_fd_sc_hd__o21ba_1 _1650_ (.A1(_0865_),
    .A2(_1031_),
    .B1_N(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__and2b_2 _1651_ (.A_N(\cpu_inst.op[0] ),
    .B(_1013_),
    .X(_1034_));
 sky130_fd_sc_hd__and3b_1 _1652_ (.A_N(\cpu_inst.op[1] ),
    .B(_1013_),
    .C(\cpu_inst.op[0] ),
    .X(_1035_));
 sky130_fd_sc_hd__nand3b_2 _1653_ (.A_N(\cpu_inst.op[1] ),
    .B(_1013_),
    .C(\cpu_inst.op[0] ),
    .Y(_1036_));
 sky130_fd_sc_hd__and2_2 _1654_ (.A(\cpu_inst.shift_right ),
    .B(_1013_),
    .X(_1037_));
 sky130_fd_sc_hd__nand2_2 _1655_ (.A(\cpu_inst.shift_right ),
    .B(_1013_),
    .Y(_1038_));
 sky130_fd_sc_hd__and2_1 _1656_ (.A(\cpu_inst.op[1] ),
    .B(_1034_),
    .X(_1039_));
 sky130_fd_sc_hd__nand2_1 _1657_ (.A(\cpu_inst.op[1] ),
    .B(_1034_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand2_1 _1658_ (.A(_1025_),
    .B(_1034_),
    .Y(_1041_));
 sky130_fd_sc_hd__mux2_1 _1659_ (.A0(_1035_),
    .A1(_1039_),
    .S(_1025_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _1660_ (.A0(_1042_),
    .A1(_1041_),
    .S(_1033_),
    .X(_1043_));
 sky130_fd_sc_hd__a221o_1 _1661_ (.A1(net76),
    .A2(_0884_),
    .B1(_1017_),
    .B2(net95),
    .C1(_0969_),
    .X(_1044_));
 sky130_fd_sc_hd__o21ba_1 _1662_ (.A1(_0873_),
    .A2(_1031_),
    .B1_N(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__inv_2 _1663_ (.A(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__mux2_1 _1664_ (.A0(_1043_),
    .A1(_1045_),
    .S(_1037_),
    .X(_1047_));
 sky130_fd_sc_hd__nor2_1 _1665_ (.A(_1027_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__a22o_1 _1666_ (.A1(\cpu_inst.PC[5] ),
    .A2(net37),
    .B1(net12),
    .B2(\cpu_inst.DI[5] ),
    .X(_1049_));
 sky130_fd_sc_hd__nor2_1 _1667_ (.A(_1015_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__xnor2_1 _1668_ (.A(net14),
    .B(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__a221o_1 _1669_ (.A1(net78),
    .A2(_0884_),
    .B1(_1017_),
    .B2(\cpu_inst.DI[5] ),
    .C1(_0961_),
    .X(_1052_));
 sky130_fd_sc_hd__a21oi_2 _1670_ (.A1(_0858_),
    .A2(_1030_),
    .B1(_1052_),
    .Y(_1053_));
 sky130_fd_sc_hd__mux2_1 _1671_ (.A0(_1040_),
    .A1(_1034_),
    .S(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nand2_1 _1672_ (.A(_1049_),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__o311a_1 _1673_ (.A1(_1035_),
    .A2(_1049_),
    .A3(_1053_),
    .B1(_1055_),
    .C1(_1038_),
    .X(_1056_));
 sky130_fd_sc_hd__a21oi_1 _1674_ (.A1(_1033_),
    .A2(_1037_),
    .B1(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__a22o_1 _1675_ (.A1(\cpu_inst.PC[4] ),
    .A2(net37),
    .B1(net12),
    .B2(\cpu_inst.DI[4] ),
    .X(_1058_));
 sky130_fd_sc_hd__or2_1 _1676_ (.A(_1015_),
    .B(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__xnor2_1 _1677_ (.A(net13),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__a2bb2o_1 _1678_ (.A1_N(_0850_),
    .A2_N(_1031_),
    .B1(_0884_),
    .B2(net79),
    .X(_0188_));
 sky130_fd_sc_hd__a211o_1 _1679_ (.A1(\cpu_inst.DI[4] ),
    .A2(_1017_),
    .B1(_0188_),
    .C1(_0957_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(_1034_),
    .A1(_1040_),
    .S(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__and3b_1 _1681_ (.A_N(_1058_),
    .B(_0189_),
    .C(_1036_),
    .X(_0191_));
 sky130_fd_sc_hd__a21oi_1 _1682_ (.A1(_1058_),
    .A2(_0190_),
    .B1(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__mux2_1 _1683_ (.A0(_1053_),
    .A1(_0192_),
    .S(_1038_),
    .X(_0193_));
 sky130_fd_sc_hd__nor2_1 _1684_ (.A(net13),
    .B(_1016_),
    .Y(_0194_));
 sky130_fd_sc_hd__a22o_1 _1685_ (.A1(\cpu_inst.PC[2] ),
    .A2(net37),
    .B1(net12),
    .B2(net98),
    .X(_0195_));
 sky130_fd_sc_hd__o21ai_1 _1686_ (.A1(net13),
    .A2(_0195_),
    .B1(_1016_),
    .Y(_0196_));
 sky130_fd_sc_hd__a21oi_1 _1687_ (.A1(net13),
    .A2(_0195_),
    .B1(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _1688_ (.A(_0194_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__a221o_1 _1689_ (.A1(net81),
    .A2(_0884_),
    .B1(_1017_),
    .B2(net98),
    .C1(_0949_),
    .X(_0199_));
 sky130_fd_sc_hd__a21o_1 _1690_ (.A1(_0834_),
    .A2(_1030_),
    .B1(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1691_ (.A0(_1034_),
    .A1(_1040_),
    .S(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__and3b_1 _1692_ (.A_N(_0195_),
    .B(_0200_),
    .C(_1036_),
    .X(_0202_));
 sky130_fd_sc_hd__a21oi_1 _1693_ (.A1(_0195_),
    .A2(_0201_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a221o_1 _1694_ (.A1(net80),
    .A2(_0884_),
    .B1(_1017_),
    .B2(net97),
    .C1(_0953_),
    .X(_0204_));
 sky130_fd_sc_hd__o21ba_1 _1695_ (.A1(_0842_),
    .A2(_1031_),
    .B1_N(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(_0203_),
    .A1(_0205_),
    .S(_1037_),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_1 _1697_ (.A1(\cpu_inst.PC[1] ),
    .A2(net37),
    .B1(net12),
    .B2(net99),
    .X(_0207_));
 sky130_fd_sc_hd__o21ai_1 _1698_ (.A1(net13),
    .A2(_0207_),
    .B1(_1016_),
    .Y(_0208_));
 sky130_fd_sc_hd__a21oi_1 _1699_ (.A1(net14),
    .A2(_0207_),
    .B1(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _1700_ (.A(_0194_),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__or2_1 _1701_ (.A(_0194_),
    .B(_0209_),
    .X(_0211_));
 sky130_fd_sc_hd__a221o_1 _1702_ (.A1(net82),
    .A2(_0884_),
    .B1(_1017_),
    .B2(net99),
    .C1(_0945_),
    .X(_0212_));
 sky130_fd_sc_hd__a21o_1 _1703_ (.A1(_0826_),
    .A2(_1030_),
    .B1(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _1704_ (.A(_1034_),
    .B(_0207_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(_1036_),
    .A1(_1040_),
    .S(_0207_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1706_ (.A0(_0214_),
    .A1(_0215_),
    .S(_0213_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1707_ (.A0(_0200_),
    .A1(_0216_),
    .S(_1038_),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _1708_ (.A1(\cpu_inst.PC[0] ),
    .A2(_0670_),
    .B1(net12),
    .B2(net100),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1709_ (.A1(net13),
    .A2(_0218_),
    .B1(_1016_),
    .Y(_0219_));
 sky130_fd_sc_hd__a21oi_1 _1710_ (.A1(net13),
    .A2(_0218_),
    .B1(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__nor2_1 _1711_ (.A(_0194_),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__or2_1 _1712_ (.A(_0194_),
    .B(_0220_),
    .X(_0222_));
 sky130_fd_sc_hd__a21o_1 _1713_ (.A1(net100),
    .A2(_1017_),
    .B1(_0940_),
    .X(_0223_));
 sky130_fd_sc_hd__a32o_1 _1714_ (.A1(_0808_),
    .A2(_0811_),
    .A3(_1030_),
    .B1(_0884_),
    .B2(net83),
    .X(_0224_));
 sky130_fd_sc_hd__o211a_1 _1715_ (.A1(_0223_),
    .A2(_0224_),
    .B1(_1039_),
    .C1(_0218_),
    .X(_0225_));
 sky130_fd_sc_hd__and2_1 _1716_ (.A(_1034_),
    .B(_0218_),
    .X(_0226_));
 sky130_fd_sc_hd__o21a_1 _1717_ (.A1(_1036_),
    .A2(_0218_),
    .B1(_1038_),
    .X(_0227_));
 sky130_fd_sc_hd__o31ai_1 _1718_ (.A1(_0223_),
    .A2(_0224_),
    .A3(_0226_),
    .B1(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__a2bb2o_1 _1719_ (.A1_N(_0225_),
    .A2_N(_0228_),
    .B1(_1037_),
    .B2(_0213_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _1720_ (.A(\cpu_inst.rotate ),
    .B(_1013_),
    .Y(_0230_));
 sky130_fd_sc_hd__o31a_1 _1721_ (.A1(\cpu_inst.load_only ),
    .A2(\cpu_inst.shift ),
    .A3(_0635_),
    .B1(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__o21ai_1 _1722_ (.A1(net42),
    .A2(_0627_),
    .B1(net84),
    .Y(_0232_));
 sky130_fd_sc_hd__and3_1 _1723_ (.A(_0574_),
    .B(_0575_),
    .C(_0641_),
    .X(_0233_));
 sky130_fd_sc_hd__nand2_1 _1724_ (.A(\cpu_inst.inc ),
    .B(_0892_),
    .Y(_0234_));
 sky130_fd_sc_hd__o2bb2a_1 _1725_ (.A1_N(\cpu_inst.compare ),
    .A2_N(_0634_),
    .B1(_0234_),
    .B2(\cpu_inst.shift ),
    .X(_0235_));
 sky130_fd_sc_hd__o221a_1 _1726_ (.A1(_0504_),
    .A2(_0231_),
    .B1(_0235_),
    .B2(\cpu_inst.rotate ),
    .C1(_0233_),
    .X(_0236_));
 sky130_fd_sc_hd__and4b_2 _1727_ (.A_N(_0590_),
    .B(_1023_),
    .C(_0232_),
    .D(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__a211oi_2 _1728_ (.A1(net13),
    .A2(_1015_),
    .B1(_1037_),
    .C1(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(_0220_),
    .A1(_0221_),
    .S(_0229_),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_1 _1730_ (.A1(_0222_),
    .A2(_0229_),
    .B1(_0238_),
    .B2(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _1731_ (.A0(_0209_),
    .A1(_0210_),
    .S(_0217_),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_1 _1732_ (.A1(_0211_),
    .A2(_0217_),
    .B1(_0240_),
    .B2(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(_0198_),
    .A1(_0197_),
    .S(_0206_),
    .X(_0243_));
 sky130_fd_sc_hd__o2bb2a_1 _1734_ (.A1_N(_0243_),
    .A2_N(_0242_),
    .B1(_0206_),
    .B2(_0198_),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _1735_ (.A1(\cpu_inst.PC[3] ),
    .A2(_0670_),
    .B1(net12),
    .B2(net97),
    .X(_0245_));
 sky130_fd_sc_hd__o21ai_1 _1736_ (.A1(net13),
    .A2(_0245_),
    .B1(_1016_),
    .Y(_0246_));
 sky130_fd_sc_hd__a21o_1 _1737_ (.A1(net13),
    .A2(_0245_),
    .B1(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2b_1 _1738_ (.A_N(_0194_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _1739_ (.A(_1034_),
    .B(_0245_),
    .Y(_0249_));
 sky130_fd_sc_hd__mux2_1 _1740_ (.A0(_1035_),
    .A1(_1039_),
    .S(_0245_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _1741_ (.A0(_0250_),
    .A1(_0249_),
    .S(_0205_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _1742_ (.A(_1038_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__o21ai_1 _1743_ (.A1(_1038_),
    .A2(_0189_),
    .B1(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__o211a_1 _1744_ (.A1(_1038_),
    .A2(_0189_),
    .B1(_0248_),
    .C1(_0252_),
    .X(_0254_));
 sky130_fd_sc_hd__a21o_1 _1745_ (.A1(_0247_),
    .A2(_0253_),
    .B1(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_1 _1746_ (.A(_0244_),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__xor2_1 _1747_ (.A(_0244_),
    .B(_0255_),
    .X(_0257_));
 sky130_fd_sc_hd__xor2_1 _1748_ (.A(_0240_),
    .B(_0241_),
    .X(_0258_));
 sky130_fd_sc_hd__xor2_1 _1749_ (.A(_0242_),
    .B(_0243_),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _1750_ (.A(_0258_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__and3_2 _1751_ (.A(\cpu_inst.adc_bcd ),
    .B(_0535_),
    .C(_0609_),
    .X(_0261_));
 sky130_fd_sc_hd__a311o_1 _1752_ (.A1(_0257_),
    .A2(_0260_),
    .A3(_0261_),
    .B1(_0256_),
    .C1(_0254_),
    .X(_0262_));
 sky130_fd_sc_hd__nor2_1 _1753_ (.A(_1015_),
    .B(_1060_),
    .Y(_0263_));
 sky130_fd_sc_hd__mux2_1 _1754_ (.A0(_1060_),
    .A1(_0263_),
    .S(_0193_),
    .X(_0264_));
 sky130_fd_sc_hd__a2bb2o_1 _1755_ (.A1_N(_1060_),
    .A2_N(_0193_),
    .B1(_0262_),
    .B2(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _1756_ (.A1(_1016_),
    .A2(_1051_),
    .B1(_1057_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21oi_1 _1757_ (.A1(_1051_),
    .A2(_1057_),
    .B1(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__a22o_1 _1758_ (.A1(_1051_),
    .A2(_1057_),
    .B1(_0265_),
    .B2(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__o21ai_1 _1759_ (.A1(_1015_),
    .A2(_1027_),
    .B1(_1047_),
    .Y(_0269_));
 sky130_fd_sc_hd__and2b_1 _1760_ (.A_N(_1048_),
    .B(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__a21oi_1 _1761_ (.A1(_0268_),
    .A2(_0269_),
    .B1(_1048_),
    .Y(_0271_));
 sky130_fd_sc_hd__a22o_1 _1762_ (.A1(\cpu_inst.PC[7] ),
    .A2(_0670_),
    .B1(_1024_),
    .B2(\cpu_inst.DI[7] ),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _1763_ (.A(_1034_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__a2bb2o_1 _1764_ (.A1_N(_1036_),
    .A2_N(_0272_),
    .B1(_0273_),
    .B2(_1045_),
    .X(_0274_));
 sky130_fd_sc_hd__a31o_1 _1765_ (.A1(_1039_),
    .A2(_1046_),
    .A3(_0272_),
    .B1(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _1766_ (.A0(_0237_),
    .A1(_0275_),
    .S(_1038_),
    .X(_0276_));
 sky130_fd_sc_hd__or2_1 _1767_ (.A(_1015_),
    .B(_0272_),
    .X(_0277_));
 sky130_fd_sc_hd__xnor2_1 _1768_ (.A(net14),
    .B(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__o21a_1 _1769_ (.A1(_1015_),
    .A2(_0278_),
    .B1(_0276_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_1 _1770_ (.A(_0276_),
    .B(_0278_),
    .Y(_0280_));
 sky130_fd_sc_hd__or2_1 _1771_ (.A(_0279_),
    .B(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__xor2_1 _1772_ (.A(_0271_),
    .B(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__xnor2_1 _1773_ (.A(_0265_),
    .B(_0267_),
    .Y(_0283_));
 sky130_fd_sc_hd__xnor2_1 _1774_ (.A(_0268_),
    .B(_0270_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand2_1 _1775_ (.A(_0283_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__a31o_1 _1776_ (.A1(_0261_),
    .A2(_0282_),
    .A3(_0285_),
    .B1(net73),
    .X(_0286_));
 sky130_fd_sc_hd__o21a_1 _1777_ (.A1(_0223_),
    .A2(_0224_),
    .B1(_1037_),
    .X(_0287_));
 sky130_fd_sc_hd__o21ba_1 _1778_ (.A1(_0271_),
    .A2(_0279_),
    .B1_N(_0280_),
    .X(_0288_));
 sky130_fd_sc_hd__xnor2_1 _1779_ (.A(_0287_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__o22a_1 _1780_ (.A1(net84),
    .A2(net63),
    .B1(_0286_),
    .B2(_0289_),
    .X(_0053_));
 sky130_fd_sc_hd__xor2_1 _1781_ (.A(_0238_),
    .B(_0239_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1782_ (.A0(net194),
    .A1(_0290_),
    .S(net65),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1783_ (.A0(\cpu_inst.ADD[1] ),
    .A1(_0258_),
    .S(net65),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(net81),
    .A1(_0259_),
    .S(net65),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1785_ (.A0(net80),
    .A1(_0257_),
    .S(net65),
    .X(_0057_));
 sky130_fd_sc_hd__xor2_1 _1786_ (.A(_0262_),
    .B(_0264_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(net79),
    .A1(_0291_),
    .S(net65),
    .X(_0058_));
 sky130_fd_sc_hd__nor2_1 _1788_ (.A(net78),
    .B(net65),
    .Y(_0292_));
 sky130_fd_sc_hd__a21oi_1 _1789_ (.A1(net65),
    .A2(_0283_),
    .B1(_0292_),
    .Y(_0059_));
 sky130_fd_sc_hd__nand2_1 _1790_ (.A(net77),
    .B(net73),
    .Y(_0293_));
 sky130_fd_sc_hd__o21ai_1 _1791_ (.A1(net73),
    .A2(_0284_),
    .B1(_0293_),
    .Y(_0060_));
 sky130_fd_sc_hd__mux2_1 _1792_ (.A0(net76),
    .A1(_0282_),
    .S(net63),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(net212),
    .A1(_0262_),
    .S(net65),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(net197),
    .A1(_1046_),
    .S(net63),
    .X(_0063_));
 sky130_fd_sc_hd__or3b_1 _1795_ (.A(net43),
    .B(_0634_),
    .C_N(_0798_),
    .X(_0294_));
 sky130_fd_sc_hd__or4b_1 _1796_ (.A(net38),
    .B(_0793_),
    .C(_0689_),
    .D_N(_0600_),
    .X(_0295_));
 sky130_fd_sc_hd__or4_1 _1797_ (.A(_0598_),
    .B(_0627_),
    .C(_0294_),
    .D(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__a32o_1 _1798_ (.A1(_0587_),
    .A2(_0675_),
    .A3(_0685_),
    .B1(_0789_),
    .B2(_0799_),
    .X(_0297_));
 sky130_fd_sc_hd__or2_1 _1799_ (.A(_0630_),
    .B(_0885_),
    .X(_0298_));
 sky130_fd_sc_hd__or4b_1 _1800_ (.A(net48),
    .B(_0296_),
    .C(net19),
    .D_N(_0297_),
    .X(_0299_));
 sky130_fd_sc_hd__or4b_1 _1801_ (.A(net94),
    .B(net87),
    .C(net50),
    .D_N(net92),
    .X(_0300_));
 sky130_fd_sc_hd__a41o_1 _1802_ (.A1(_0639_),
    .A2(_0682_),
    .A3(_0730_),
    .A4(_0300_),
    .B1(_0602_),
    .X(_0301_));
 sky130_fd_sc_hd__or4b_1 _1803_ (.A(net46),
    .B(_0882_),
    .C(_1022_),
    .D_N(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__nor3_1 _1804_ (.A(_1019_),
    .B(_0299_),
    .C(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__nor3_2 _1805_ (.A(_0755_),
    .B(_1028_),
    .C(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__mux2_1 _1806_ (.A0(net230),
    .A1(_0943_),
    .S(net5),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(net246),
    .A1(_0947_),
    .S(net5),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1808_ (.A0(net234),
    .A1(_0951_),
    .S(net6),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1809_ (.A0(net233),
    .A1(_0955_),
    .S(net5),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(net240),
    .A1(_0959_),
    .S(net5),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1811_ (.A0(net236),
    .A1(_0963_),
    .S(net5),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1812_ (.A0(net229),
    .A1(_0967_),
    .S(net5),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(net235),
    .A1(_0971_),
    .S(net5),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1814_ (.A0(net214),
    .A1(_0902_),
    .S(net5),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1815_ (.A0(net213),
    .A1(_0907_),
    .S(net5),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1816_ (.A0(net218),
    .A1(_0912_),
    .S(net5),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1817_ (.A0(net227),
    .A1(_0917_),
    .S(net6),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1818_ (.A0(net220),
    .A1(_0922_),
    .S(net6),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(net204),
    .A1(_0927_),
    .S(net6),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1820_ (.A0(net206),
    .A1(_0932_),
    .S(net6),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1821_ (.A0(net216),
    .A1(_0937_),
    .S(net6),
    .X(_0079_));
 sky130_fd_sc_hd__and3_1 _1822_ (.A(\cpu_inst.D ),
    .B(\cpu_inst.adc_sbc ),
    .C(net63),
    .X(_0305_));
 sky130_fd_sc_hd__a21o_1 _1823_ (.A1(net242),
    .A2(net73),
    .B1(_0305_),
    .X(_0080_));
 sky130_fd_sc_hd__a2bb2o_1 _1824_ (.A1_N(\cpu_inst.write_back ),
    .A2_N(net47),
    .B1(_0632_),
    .B2(\cpu_inst.shift ),
    .X(_0306_));
 sky130_fd_sc_hd__or3_1 _1825_ (.A(\cpu_inst.compare ),
    .B(\cpu_inst.shift ),
    .C(\cpu_inst.adc_sbc ),
    .X(_0307_));
 sky130_fd_sc_hd__or4_1 _1826_ (.A(net74),
    .B(\cpu_inst.clc ),
    .C(\cpu_inst.sec ),
    .D(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__or3_1 _1827_ (.A(\cpu_inst.write_back ),
    .B(net47),
    .C(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__o211a_1 _1828_ (.A1(_0554_),
    .A2(_0306_),
    .B1(_0309_),
    .C1(net60),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(_0505_),
    .A1(net83),
    .S(net74),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(_0311_),
    .A1(net84),
    .S(_0307_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _1831_ (.A0(net100),
    .A1(_0312_),
    .S(_0555_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(\cpu_inst.C ),
    .A1(_0313_),
    .S(_0310_),
    .X(_0081_));
 sky130_fd_sc_hd__or2_1 _1833_ (.A(_0539_),
    .B(net38),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _1834_ (.A(net27),
    .B(_0758_),
    .Y(_0315_));
 sky130_fd_sc_hd__o21a_1 _1835_ (.A1(_0554_),
    .A2(_0314_),
    .B1(net60),
    .X(_0316_));
 sky130_fd_sc_hd__a2111o_1 _1836_ (.A1(\cpu_inst.load_reg ),
    .A2(_0809_),
    .B1(\cpu_inst.compare ),
    .C1(net74),
    .D1(net47),
    .X(_0317_));
 sky130_fd_sc_hd__o21a_1 _1837_ (.A1(\cpu_inst.bit_ins ),
    .A2(_0317_),
    .B1(_0316_),
    .X(_0318_));
 sky130_fd_sc_hd__o21ba_1 _1838_ (.A1(net74),
    .A2(_0554_),
    .B1_N(net38),
    .X(_0319_));
 sky130_fd_sc_hd__or4_1 _1839_ (.A(net81),
    .B(net82),
    .C(net83),
    .D(net76),
    .X(_0320_));
 sky130_fd_sc_hd__or4_1 _1840_ (.A(net78),
    .B(net77),
    .C(net79),
    .D(net80),
    .X(_0321_));
 sky130_fd_sc_hd__nor2_1 _1841_ (.A(_0320_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__mux2_1 _1842_ (.A0(net99),
    .A1(net82),
    .S(_0555_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _1843_ (.A0(_0322_),
    .A1(_0323_),
    .S(_0319_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(net238),
    .A1(_0324_),
    .S(_0318_),
    .X(_0082_));
 sky130_fd_sc_hd__a31o_1 _1845_ (.A1(\cpu_inst.bit_ins ),
    .A2(net60),
    .A3(_0634_),
    .B1(_0315_),
    .X(_0325_));
 sky130_fd_sc_hd__a31o_1 _1846_ (.A1(\cpu_inst.bit_ins ),
    .A2(net60),
    .A3(_0634_),
    .B1(_0316_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _1847_ (.A(_0317_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__mux2_1 _1848_ (.A0(net95),
    .A1(net76),
    .S(_0314_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _1849_ (.A0(_0328_),
    .A1(net222),
    .S(_0327_),
    .X(_0083_));
 sky130_fd_sc_hd__o41a_1 _1850_ (.A1(net74),
    .A2(\cpu_inst.cld ),
    .A3(\cpu_inst.sed ),
    .A4(net47),
    .B1(_0315_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _1851_ (.A0(_0507_),
    .A1(net80),
    .S(net74),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _1852_ (.A0(net97),
    .A1(_0330_),
    .S(_0555_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _1853_ (.A0(\cpu_inst.D ),
    .A1(_0331_),
    .S(_0329_),
    .X(_0084_));
 sky130_fd_sc_hd__or4_1 _1854_ (.A(net48),
    .B(_0554_),
    .C(_0568_),
    .D(_0729_),
    .X(_0332_));
 sky130_fd_sc_hd__o21a_1 _1855_ (.A1(net74),
    .A2(_0526_),
    .B1(net59),
    .X(_0333_));
 sky130_fd_sc_hd__o311a_1 _1856_ (.A1(\cpu_inst.cli ),
    .A2(\cpu_inst.sei ),
    .A3(_0730_),
    .B1(_0332_),
    .C1(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _1857_ (.A0(_0501_),
    .A1(\cpu_inst.cli ),
    .S(_0729_),
    .X(_0335_));
 sky130_fd_sc_hd__nor2_1 _1858_ (.A(_0554_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__a211o_1 _1859_ (.A1(net98),
    .A2(_0554_),
    .B1(_0568_),
    .C1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(net254),
    .A1(_0337_),
    .S(_0334_),
    .X(_0085_));
 sky130_fd_sc_hd__o41a_1 _1861_ (.A1(net74),
    .A2(\cpu_inst.clv ),
    .A3(\cpu_inst.adc_sbc ),
    .A4(net47),
    .B1(_0325_),
    .X(_0338_));
 sky130_fd_sc_hd__xnor2_1 _1862_ (.A(\cpu_inst.ALU.BI7 ),
    .B(\cpu_inst.ALU.AI7 ),
    .Y(_0339_));
 sky130_fd_sc_hd__xnor2_1 _1863_ (.A(\cpu_inst.ALU.CO ),
    .B(net76),
    .Y(_0340_));
 sky130_fd_sc_hd__a211oi_1 _1864_ (.A1(_0339_),
    .A2(_0340_),
    .B1(net74),
    .C1(\cpu_inst.clv ),
    .Y(_0341_));
 sky130_fd_sc_hd__o21ai_1 _1865_ (.A1(_0339_),
    .A2(_0340_),
    .B1(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__a21oi_1 _1866_ (.A1(\cpu_inst.plp ),
    .A2(net77),
    .B1(_0540_),
    .Y(_0343_));
 sky130_fd_sc_hd__o2bb2a_1 _1867_ (.A1_N(_0342_),
    .A2_N(_0343_),
    .B1(net96),
    .B2(net48),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _1868_ (.A0(net217),
    .A1(_0344_),
    .S(_0338_),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _1869_ (.A1(net75),
    .A2(net26),
    .B1(_1028_),
    .B2(net59),
    .X(_0087_));
 sky130_fd_sc_hd__and3_2 _1870_ (.A(net102),
    .B(net59),
    .C(_1028_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _1871_ (.A0(net154),
    .A1(net100),
    .S(_0345_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1872_ (.A0(net140),
    .A1(net99),
    .S(_0345_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1873_ (.A0(net173),
    .A1(net98),
    .S(_0345_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1874_ (.A0(net149),
    .A1(net97),
    .S(_0345_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1875_ (.A0(net161),
    .A1(\cpu_inst.DI[4] ),
    .S(_0345_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1876_ (.A0(net237),
    .A1(\cpu_inst.DI[5] ),
    .S(_0345_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1877_ (.A0(net153),
    .A1(net96),
    .S(_0345_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _1878_ (.A0(net164),
    .A1(net95),
    .S(_0345_),
    .X(_0095_));
 sky130_fd_sc_hd__nor2_1 _1879_ (.A(_0510_),
    .B(_0539_),
    .Y(_0096_));
 sky130_fd_sc_hd__or2_2 _1880_ (.A(_0622_),
    .B(_0648_),
    .X(_0346_));
 sky130_fd_sc_hd__nor2_2 _1881_ (.A(_0655_),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__nor2_1 _1882_ (.A(_0613_),
    .B(_0732_),
    .Y(_0348_));
 sky130_fd_sc_hd__or2_1 _1883_ (.A(_0613_),
    .B(_0732_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _1884_ (.A(_0531_),
    .B(_0656_),
    .Y(_0350_));
 sky130_fd_sc_hd__nor2_1 _1885_ (.A(_0654_),
    .B(_0346_),
    .Y(_0351_));
 sky130_fd_sc_hd__or3_1 _1886_ (.A(_0614_),
    .B(_0346_),
    .C(_0350_),
    .X(_0352_));
 sky130_fd_sc_hd__a21bo_1 _1887_ (.A1(_0347_),
    .A2(_0348_),
    .B1_N(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__a21oi_1 _1888_ (.A1(_0620_),
    .A2(_0654_),
    .B1(_0617_),
    .Y(_0354_));
 sky130_fd_sc_hd__a31o_1 _1889_ (.A1(_0546_),
    .A2(_0622_),
    .A3(_0348_),
    .B1(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__and3_1 _1890_ (.A(_0543_),
    .B(_0348_),
    .C(_0351_),
    .X(_0356_));
 sky130_fd_sc_hd__o21a_1 _1891_ (.A1(_0546_),
    .A2(_0347_),
    .B1(_0664_),
    .X(_0357_));
 sky130_fd_sc_hd__and3_2 _1892_ (.A(_0530_),
    .B(_0620_),
    .C(_0648_),
    .X(_0358_));
 sky130_fd_sc_hd__or3b_1 _1893_ (.A(_0545_),
    .B(_0656_),
    .C_N(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _1894_ (.A(_0349_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__nand2_1 _1895_ (.A(net29),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__a211o_1 _1896_ (.A1(_0619_),
    .A2(_0349_),
    .B1(_0346_),
    .C1(_0697_),
    .X(_0362_));
 sky130_fd_sc_hd__or4b_1 _1897_ (.A(_0356_),
    .B(_0357_),
    .C(_0361_),
    .D_N(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_1 _1898_ (.A(_0546_),
    .B(_0665_),
    .Y(_0364_));
 sky130_fd_sc_hd__or2_1 _1899_ (.A(net28),
    .B(_0356_),
    .X(_0365_));
 sky130_fd_sc_hd__o32a_1 _1900_ (.A1(_0353_),
    .A2(_0355_),
    .A3(_0363_),
    .B1(net30),
    .B2(net248),
    .X(_0097_));
 sky130_fd_sc_hd__a211oi_2 _1901_ (.A1(_0697_),
    .A2(_0350_),
    .B1(_0346_),
    .C1(_0644_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(net30),
    .B(_0666_),
    .Y(_0367_));
 sky130_fd_sc_hd__o22a_1 _1903_ (.A1(\cpu_inst.dst_reg[0] ),
    .A2(net30),
    .B1(_0366_),
    .B2(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__a31o_1 _1904_ (.A1(_0671_),
    .A2(_0347_),
    .A3(_0348_),
    .B1(_0368_),
    .X(_0098_));
 sky130_fd_sc_hd__nor2_1 _1905_ (.A(_0622_),
    .B(_0666_),
    .Y(_0369_));
 sky130_fd_sc_hd__and3_1 _1906_ (.A(_0544_),
    .B(_0664_),
    .C(_0358_),
    .X(_0370_));
 sky130_fd_sc_hd__a211o_1 _1907_ (.A1(_0731_),
    .A2(_0351_),
    .B1(_0366_),
    .C1(_0369_),
    .X(_0371_));
 sky130_fd_sc_hd__o32a_1 _1908_ (.A1(_0361_),
    .A2(_0370_),
    .A3(_0371_),
    .B1(net29),
    .B2(net136),
    .X(_0099_));
 sky130_fd_sc_hd__and2b_1 _1909_ (.A_N(_0648_),
    .B(_0369_),
    .X(_0372_));
 sky130_fd_sc_hd__nand2_1 _1910_ (.A(_0531_),
    .B(_0347_),
    .Y(_0373_));
 sky130_fd_sc_hd__a21oi_1 _1911_ (.A1(_0359_),
    .A2(_0373_),
    .B1(_0644_),
    .Y(_0374_));
 sky130_fd_sc_hd__a211o_1 _1912_ (.A1(_0347_),
    .A2(_0364_),
    .B1(_0372_),
    .C1(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__o22a_1 _1913_ (.A1(net196),
    .A2(net29),
    .B1(_0365_),
    .B2(_0375_),
    .X(_0100_));
 sky130_fd_sc_hd__nor2_1 _1914_ (.A(_0614_),
    .B(_0373_),
    .Y(_0376_));
 sky130_fd_sc_hd__a221o_1 _1915_ (.A1(_0347_),
    .A2(_0348_),
    .B1(_0358_),
    .B2(_0698_),
    .C1(_0361_),
    .X(_0377_));
 sky130_fd_sc_hd__o32a_1 _1916_ (.A1(_0375_),
    .A2(_0376_),
    .A3(_0377_),
    .B1(net29),
    .B2(\cpu_inst.src_reg[1] ),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _1917_ (.A(_0531_),
    .B(_0731_),
    .X(_0378_));
 sky130_fd_sc_hd__or3b_1 _1918_ (.A(_0544_),
    .B(_0346_),
    .C_N(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__o221a_1 _1919_ (.A1(_0613_),
    .A2(_0617_),
    .B1(_0693_),
    .B2(_0546_),
    .C1(net30),
    .X(_0380_));
 sky130_fd_sc_hd__o2bb2a_1 _1920_ (.A1_N(_0379_),
    .A2_N(_0380_),
    .B1(net195),
    .B2(net29),
    .X(_0102_));
 sky130_fd_sc_hd__a21o_1 _1921_ (.A1(_0618_),
    .A2(_0347_),
    .B1(net28),
    .X(_0381_));
 sky130_fd_sc_hd__o22a_1 _1922_ (.A1(\cpu_inst.store ),
    .A2(net29),
    .B1(_0376_),
    .B2(_0381_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _1923_ (.A(\cpu_inst.write_back ),
    .B(net28),
    .X(_0382_));
 sky130_fd_sc_hd__a31o_1 _1924_ (.A1(net29),
    .A2(_0346_),
    .A3(_0378_),
    .B1(_0382_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1925_ (.A0(net243),
    .A1(_0351_),
    .S(net31),
    .X(_0105_));
 sky130_fd_sc_hd__a31o_1 _1926_ (.A1(_0656_),
    .A2(_0358_),
    .A3(_0378_),
    .B1(_0370_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _1927_ (.A0(net198),
    .A1(_0383_),
    .S(net29),
    .X(_0106_));
 sky130_fd_sc_hd__o21a_1 _1928_ (.A1(net48),
    .A2(_0686_),
    .B1(net59),
    .X(_0384_));
 sky130_fd_sc_hd__nor2_1 _1929_ (.A(_0649_),
    .B(_0654_),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _1930_ (.A(_0618_),
    .B(_0650_),
    .C(_0655_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _1931_ (.A0(\cpu_inst.adc_sbc ),
    .A1(_0386_),
    .S(_0384_),
    .X(_0107_));
 sky130_fd_sc_hd__and3b_1 _1932_ (.A_N(_0667_),
    .B(_0731_),
    .C(_0645_),
    .X(_0387_));
 sky130_fd_sc_hd__a21o_1 _1933_ (.A1(net244),
    .A2(net27),
    .B1(_0387_),
    .X(_0108_));
 sky130_fd_sc_hd__and3_1 _1934_ (.A(\cpu_inst.D ),
    .B(_0622_),
    .C(_0386_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _1935_ (.A0(\cpu_inst.adc_bcd ),
    .A1(_0388_),
    .S(_0384_),
    .X(_0109_));
 sky130_fd_sc_hd__or3_1 _1936_ (.A(_0545_),
    .B(_0612_),
    .C(_0644_),
    .X(_0389_));
 sky130_fd_sc_hd__o211a_1 _1937_ (.A1(_0617_),
    .A2(_0655_),
    .B1(_0762_),
    .C1(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__and2b_1 _1938_ (.A_N(_0390_),
    .B(_0358_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _1939_ (.A0(net257),
    .A1(_0391_),
    .S(_0541_),
    .X(_0110_));
 sky130_fd_sc_hd__and2_1 _1940_ (.A(\cpu_inst.shift_right ),
    .B(net27),
    .X(_0392_));
 sky130_fd_sc_hd__a31o_1 _1941_ (.A1(net31),
    .A2(_0651_),
    .A3(_0731_),
    .B1(_0392_),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _1942_ (.A1(net228),
    .A2(net27),
    .B1(_0656_),
    .B2(_0387_),
    .X(_0112_));
 sky130_fd_sc_hd__or2_1 _1943_ (.A(\cpu_inst.op[0] ),
    .B(net31),
    .X(_0393_));
 sky130_fd_sc_hd__or3_1 _1944_ (.A(_0617_),
    .B(_0621_),
    .C(_0385_),
    .X(_0394_));
 sky130_fd_sc_hd__o31a_1 _1945_ (.A1(net27),
    .A2(_0656_),
    .A3(_0394_),
    .B1(_0393_),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _1946_ (.A1(_0651_),
    .A2(_0731_),
    .B1(_0358_),
    .B2(_0618_),
    .X(_0395_));
 sky130_fd_sc_hd__nor3_1 _1947_ (.A(_0644_),
    .B(_0715_),
    .C(_0350_),
    .Y(_0396_));
 sky130_fd_sc_hd__or4bb_1 _1948_ (.A(_0395_),
    .B(net11),
    .C_N(_0360_),
    .D_N(_0394_),
    .X(_0397_));
 sky130_fd_sc_hd__a31o_1 _1949_ (.A1(_0654_),
    .A2(_0358_),
    .A3(_0378_),
    .B1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__or3_1 _1950_ (.A(_0372_),
    .B(_0391_),
    .C(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _1951_ (.A(net31),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__o32a_1 _1952_ (.A1(_0713_),
    .A2(_0731_),
    .A3(_0400_),
    .B1(net31),
    .B2(\cpu_inst.op[1] ),
    .X(_0114_));
 sky130_fd_sc_hd__a21bo_1 _1953_ (.A1(net150),
    .A2(net27),
    .B1_N(_0400_),
    .X(_0115_));
 sky130_fd_sc_hd__a21o_1 _1954_ (.A1(_0714_),
    .A2(_0731_),
    .B1(_0399_),
    .X(_0401_));
 sky130_fd_sc_hd__nor2_1 _1955_ (.A(net26),
    .B(_0620_),
    .Y(_0402_));
 sky130_fd_sc_hd__a22o_1 _1956_ (.A1(\cpu_inst.op[3] ),
    .A2(net26),
    .B1(_0401_),
    .B2(_0402_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1957_ (.A0(net250),
    .A1(net11),
    .S(net31),
    .X(_0117_));
 sky130_fd_sc_hd__and3_1 _1958_ (.A(net31),
    .B(_0543_),
    .C(_0664_),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _1959_ (.A1(net247),
    .A2(net26),
    .B1(_0351_),
    .B2(_0403_),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _1960_ (.A(\cpu_inst.sei ),
    .B(net26),
    .X(_0404_));
 sky130_fd_sc_hd__a31o_1 _1961_ (.A1(_0364_),
    .A2(_0385_),
    .A3(_0402_),
    .B1(_0404_),
    .X(_0119_));
 sky130_fd_sc_hd__and3_1 _1962_ (.A(net31),
    .B(_0654_),
    .C(_0364_),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _1963_ (.A1(net239),
    .A2(net26),
    .B1(_0651_),
    .B2(_0405_),
    .X(_0120_));
 sky130_fd_sc_hd__and3_1 _1964_ (.A(net31),
    .B(_0545_),
    .C(_0655_),
    .X(_0406_));
 sky130_fd_sc_hd__a32o_1 _1965_ (.A1(_0664_),
    .A2(_0358_),
    .A3(_0406_),
    .B1(net26),
    .B2(net190),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _1966_ (.A1(net277),
    .A2(net26),
    .B1(_0358_),
    .B2(_0405_),
    .X(_0122_));
 sky130_fd_sc_hd__a32o_1 _1967_ (.A1(_0664_),
    .A2(_0714_),
    .A3(_0406_),
    .B1(net26),
    .B2(net138),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _1968_ (.A1(net231),
    .A2(net26),
    .B1(_0714_),
    .B2(_0405_),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _1969_ (.A1(\cpu_inst.php ),
    .A2(net27),
    .B1(_0649_),
    .B2(_0668_),
    .X(_0125_));
 sky130_fd_sc_hd__nor2_1 _1970_ (.A(_0665_),
    .B(_0715_),
    .Y(_0407_));
 sky130_fd_sc_hd__mux2_1 _1971_ (.A0(\cpu_inst.plp ),
    .A1(_0407_),
    .S(net29),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1972_ (.A0(net202),
    .A1(_0656_),
    .S(net56),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1973_ (.A0(net225),
    .A1(_0650_),
    .S(net59),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1974_ (.A0(net200),
    .A1(_0621_),
    .S(net59),
    .X(_0129_));
 sky130_fd_sc_hd__o221a_1 _1975_ (.A1(net53),
    .A2(_0675_),
    .B1(_0680_),
    .B2(_0602_),
    .C1(_0633_),
    .X(_0408_));
 sky130_fd_sc_hd__a2111oi_1 _1976_ (.A1(net49),
    .A2(net48),
    .B1(_0568_),
    .C1(_0588_),
    .D1(net37),
    .Y(_0409_));
 sky130_fd_sc_hd__and3_2 _1977_ (.A(_0739_),
    .B(_0408_),
    .C(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__or4b_1 _1978_ (.A(_0539_),
    .B(net19),
    .C(net43),
    .D_N(_1018_),
    .X(_0411_));
 sky130_fd_sc_hd__a21bo_2 _1979_ (.A1(_0530_),
    .A2(net48),
    .B1_N(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__or2_2 _1980_ (.A(net43),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_1 _1981_ (.A(_0530_),
    .B(_0540_),
    .Y(_0414_));
 sky130_fd_sc_hd__a221o_1 _1982_ (.A1(net83),
    .A2(net18),
    .B1(net21),
    .B2(\cpu_inst.ABL[0] ),
    .C1(_0899_),
    .X(_0415_));
 sky130_fd_sc_hd__a21o_1 _1983_ (.A1(\cpu_inst.PC[0] ),
    .A2(_0413_),
    .B1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__nand2b_1 _1984_ (.A_N(_0410_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__xnor2_1 _1985_ (.A(_0410_),
    .B(_0416_),
    .Y(_0418_));
 sky130_fd_sc_hd__mux2_1 _1986_ (.A0(\cpu_inst.PC[0] ),
    .A1(_0418_),
    .S(net65),
    .X(_0130_));
 sky130_fd_sc_hd__o21a_1 _1987_ (.A1(net40),
    .A2(net19),
    .B1(\cpu_inst.ADD[1] ),
    .X(_0419_));
 sky130_fd_sc_hd__a221o_1 _1988_ (.A1(_0510_),
    .A2(_0566_),
    .B1(net22),
    .B2(\cpu_inst.ABL[1] ),
    .C1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__a21oi_1 _1989_ (.A1(\cpu_inst.PC[1] ),
    .A2(_0413_),
    .B1(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__or2_1 _1990_ (.A(_0417_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _1991_ (.A(_0417_),
    .B(_0421_),
    .Y(_0423_));
 sky130_fd_sc_hd__and2_1 _1992_ (.A(\cpu_inst.PC[1] ),
    .B(net73),
    .X(_0424_));
 sky130_fd_sc_hd__a31o_1 _1993_ (.A1(net64),
    .A2(_0422_),
    .A3(_0423_),
    .B1(_0424_),
    .X(_0131_));
 sky130_fd_sc_hd__o21a_1 _1994_ (.A1(_0499_),
    .A2(\cpu_inst.res ),
    .B1(net46),
    .X(_0425_));
 sky130_fd_sc_hd__a221o_1 _1995_ (.A1(net81),
    .A2(net40),
    .B1(net21),
    .B2(\cpu_inst.ABL[2] ),
    .C1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__a221o_1 _1996_ (.A1(\cpu_inst.ADD[2] ),
    .A2(net18),
    .B1(_0413_),
    .B2(\cpu_inst.PC[2] ),
    .C1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__and2b_1 _1997_ (.A_N(_0422_),
    .B(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__and2b_1 _1998_ (.A_N(_0427_),
    .B(_0422_),
    .X(_0429_));
 sky130_fd_sc_hd__nor2_1 _1999_ (.A(_0428_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__mux2_1 _2000_ (.A0(\cpu_inst.PC[2] ),
    .A1(_0430_),
    .S(net66),
    .X(_0132_));
 sky130_fd_sc_hd__a221o_1 _2001_ (.A1(net80),
    .A2(net40),
    .B1(net22),
    .B2(\cpu_inst.ABL[3] ),
    .C1(_0566_),
    .X(_0431_));
 sky130_fd_sc_hd__a221o_1 _2002_ (.A1(\cpu_inst.ADD[3] ),
    .A2(net18),
    .B1(_0413_),
    .B2(\cpu_inst.PC[3] ),
    .C1(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__xor2_1 _2003_ (.A(_0428_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _2004_ (.A0(\cpu_inst.PC[3] ),
    .A1(_0433_),
    .S(net64),
    .X(_0133_));
 sky130_fd_sc_hd__a221o_1 _2005_ (.A1(net79),
    .A2(net40),
    .B1(net22),
    .B2(\cpu_inst.ABL[4] ),
    .C1(net46),
    .X(_0434_));
 sky130_fd_sc_hd__a221o_1 _2006_ (.A1(net79),
    .A2(net18),
    .B1(_0413_),
    .B2(\cpu_inst.PC[4] ),
    .C1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__and3_1 _2007_ (.A(_0428_),
    .B(_0432_),
    .C(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__a21oi_1 _2008_ (.A1(_0428_),
    .A2(_0432_),
    .B1(_0435_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _2009_ (.A(net241),
    .B(net73),
    .Y(_0438_));
 sky130_fd_sc_hd__o31ai_1 _2010_ (.A1(net73),
    .A2(_0436_),
    .A3(_0437_),
    .B1(_0438_),
    .Y(_0134_));
 sky130_fd_sc_hd__a221o_1 _2011_ (.A1(\cpu_inst.ADD[5] ),
    .A2(net40),
    .B1(net22),
    .B2(\cpu_inst.ABL[5] ),
    .C1(_0566_),
    .X(_0439_));
 sky130_fd_sc_hd__a221o_1 _2012_ (.A1(\cpu_inst.ADD[5] ),
    .A2(net18),
    .B1(_0413_),
    .B2(\cpu_inst.PC[5] ),
    .C1(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__nor2_1 _2013_ (.A(_0436_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__and2_1 _2014_ (.A(_0436_),
    .B(_0440_),
    .X(_0442_));
 sky130_fd_sc_hd__nor2_1 _2015_ (.A(_0441_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__mux2_1 _2016_ (.A0(\cpu_inst.PC[5] ),
    .A1(_0443_),
    .S(net66),
    .X(_0135_));
 sky130_fd_sc_hd__a221o_1 _2017_ (.A1(\cpu_inst.ADD[6] ),
    .A2(net39),
    .B1(net22),
    .B2(\cpu_inst.ABL[6] ),
    .C1(net45),
    .X(_0444_));
 sky130_fd_sc_hd__a221o_1 _2018_ (.A1(net77),
    .A2(net18),
    .B1(_0413_),
    .B2(\cpu_inst.PC[6] ),
    .C1(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__and3_1 _2019_ (.A(_0436_),
    .B(_0440_),
    .C(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__nor2_1 _2020_ (.A(_0442_),
    .B(_0445_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _2021_ (.A(_0446_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__mux2_1 _2022_ (.A0(\cpu_inst.PC[6] ),
    .A1(_0448_),
    .S(net66),
    .X(_0136_));
 sky130_fd_sc_hd__a221o_1 _2023_ (.A1(net76),
    .A2(net39),
    .B1(net22),
    .B2(\cpu_inst.ABL[7] ),
    .C1(net45),
    .X(_0449_));
 sky130_fd_sc_hd__a221o_1 _2024_ (.A1(\cpu_inst.ADD[7] ),
    .A2(net18),
    .B1(_0413_),
    .B2(\cpu_inst.PC[7] ),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__xor2_1 _2025_ (.A(_0446_),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _2026_ (.A0(\cpu_inst.PC[7] ),
    .A1(_0451_),
    .S(net64),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _2027_ (.A1(net83),
    .A2(net43),
    .B1(net21),
    .B2(\cpu_inst.ABH[0] ),
    .X(_0452_));
 sky130_fd_sc_hd__or3_1 _2028_ (.A(net45),
    .B(_0940_),
    .C(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__a221o_1 _2029_ (.A1(net100),
    .A2(net18),
    .B1(_0412_),
    .B2(\cpu_inst.PC[8] ),
    .C1(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__and3_1 _2030_ (.A(_0446_),
    .B(_0450_),
    .C(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__a21oi_1 _2031_ (.A1(_0446_),
    .A2(_0450_),
    .B1(_0454_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _2032_ (.A(net224),
    .B(net73),
    .Y(_0457_));
 sky130_fd_sc_hd__o31ai_1 _2033_ (.A1(net73),
    .A2(_0455_),
    .A3(_0456_),
    .B1(_0457_),
    .Y(_0138_));
 sky130_fd_sc_hd__a22o_1 _2034_ (.A1(net82),
    .A2(net43),
    .B1(net21),
    .B2(\cpu_inst.ABH[1] ),
    .X(_0458_));
 sky130_fd_sc_hd__or3_1 _2035_ (.A(net45),
    .B(_0945_),
    .C(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__a221o_1 _2036_ (.A1(net99),
    .A2(net18),
    .B1(_0412_),
    .B2(\cpu_inst.PC[9] ),
    .C1(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__xor2_1 _2037_ (.A(_0455_),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _2038_ (.A0(net274),
    .A1(_0461_),
    .S(net66),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_1 _2039_ (.A1(net81),
    .A2(net43),
    .B1(net21),
    .B2(\cpu_inst.ABH[2] ),
    .X(_0462_));
 sky130_fd_sc_hd__or3_1 _2040_ (.A(net45),
    .B(_0949_),
    .C(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__a221o_1 _2041_ (.A1(net98),
    .A2(net18),
    .B1(_0412_),
    .B2(\cpu_inst.PC[10] ),
    .C1(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__and3_1 _2042_ (.A(_0455_),
    .B(_0460_),
    .C(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__a21oi_1 _2043_ (.A1(_0455_),
    .A2(_0460_),
    .B1(_0464_),
    .Y(_0466_));
 sky130_fd_sc_hd__nor2_1 _2044_ (.A(_0465_),
    .B(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__mux2_1 _2045_ (.A0(net270),
    .A1(_0467_),
    .S(net62),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _2046_ (.A1(net80),
    .A2(_0578_),
    .B1(net21),
    .B2(\cpu_inst.ABH[3] ),
    .X(_0468_));
 sky130_fd_sc_hd__or3_1 _2047_ (.A(net45),
    .B(_0953_),
    .C(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a221o_1 _2048_ (.A1(net97),
    .A2(net19),
    .B1(_0412_),
    .B2(\cpu_inst.PC[11] ),
    .C1(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__xor2_1 _2049_ (.A(_0465_),
    .B(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _2050_ (.A0(net253),
    .A1(_0471_),
    .S(net62),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_1 _2051_ (.A1(net79),
    .A2(_0578_),
    .B1(net21),
    .B2(\cpu_inst.ABH[4] ),
    .X(_0472_));
 sky130_fd_sc_hd__or3_1 _2052_ (.A(net45),
    .B(_0957_),
    .C(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__a221o_1 _2053_ (.A1(\cpu_inst.DI[4] ),
    .A2(net19),
    .B1(_0412_),
    .B2(\cpu_inst.PC[12] ),
    .C1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__and3_1 _2054_ (.A(_0465_),
    .B(_0470_),
    .C(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__a21oi_1 _2055_ (.A1(_0465_),
    .A2(_0470_),
    .B1(_0474_),
    .Y(_0476_));
 sky130_fd_sc_hd__nor2_1 _2056_ (.A(_0475_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__mux2_1 _2057_ (.A0(net279),
    .A1(_0477_),
    .S(net62),
    .X(_0142_));
 sky130_fd_sc_hd__a22o_1 _2058_ (.A1(net78),
    .A2(_0578_),
    .B1(net21),
    .B2(\cpu_inst.ABH[5] ),
    .X(_0478_));
 sky130_fd_sc_hd__or3_1 _2059_ (.A(net45),
    .B(_0961_),
    .C(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__a221o_1 _2060_ (.A1(\cpu_inst.DI[5] ),
    .A2(net19),
    .B1(_0412_),
    .B2(\cpu_inst.PC[13] ),
    .C1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__nor2_1 _2061_ (.A(_0475_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__and2_1 _2062_ (.A(_0475_),
    .B(_0480_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _2063_ (.A(net211),
    .B(net72),
    .Y(_0483_));
 sky130_fd_sc_hd__o31ai_1 _2064_ (.A1(net72),
    .A2(_0481_),
    .A3(_0482_),
    .B1(_0483_),
    .Y(_0143_));
 sky130_fd_sc_hd__a22o_1 _2065_ (.A1(net77),
    .A2(net43),
    .B1(net21),
    .B2(\cpu_inst.ABH[6] ),
    .X(_0484_));
 sky130_fd_sc_hd__or3_1 _2066_ (.A(net46),
    .B(_0965_),
    .C(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__a221o_1 _2067_ (.A1(net96),
    .A2(net19),
    .B1(_0412_),
    .B2(\cpu_inst.PC[14] ),
    .C1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__nand2_1 _2068_ (.A(_0482_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__or2_1 _2069_ (.A(_0482_),
    .B(_0486_),
    .X(_0488_));
 sky130_fd_sc_hd__and2_1 _2070_ (.A(\cpu_inst.PC[14] ),
    .B(net71),
    .X(_0489_));
 sky130_fd_sc_hd__a31o_1 _2071_ (.A1(net61),
    .A2(_0487_),
    .A3(_0488_),
    .B1(_0489_),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_1 _2072_ (.A1(net76),
    .A2(net43),
    .B1(net21),
    .B2(\cpu_inst.ABH[7] ),
    .X(_0490_));
 sky130_fd_sc_hd__or3_1 _2073_ (.A(net46),
    .B(_0969_),
    .C(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__a221o_1 _2074_ (.A1(net95),
    .A2(net19),
    .B1(_0412_),
    .B2(\cpu_inst.PC[15] ),
    .C1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__xnor2_1 _2075_ (.A(_0487_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__mux2_1 _2076_ (.A0(net269),
    .A1(_0493_),
    .S(net61),
    .X(_0145_));
 sky130_fd_sc_hd__a21oi_1 _2077_ (.A1(net60),
    .A2(_0568_),
    .B1(_0499_),
    .Y(_0494_));
 sky130_fd_sc_hd__a31o_1 _2078_ (.A1(_0499_),
    .A2(net3),
    .A3(_0509_),
    .B1(_0494_),
    .X(_0146_));
 sky130_fd_sc_hd__nor3_1 _2079_ (.A(net16),
    .B(_0805_),
    .C(_0977_),
    .Y(_0495_));
 sky130_fd_sc_hd__mux2_1 _2080_ (.A0(net199),
    .A1(_0980_),
    .S(_0495_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2081_ (.A0(net144),
    .A1(_0987_),
    .S(net10),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2082_ (.A0(net143),
    .A1(_0992_),
    .S(net10),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2083_ (.A0(net137),
    .A1(_0996_),
    .S(net10),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2084_ (.A0(net135),
    .A1(_0997_),
    .S(net10),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2085_ (.A0(net142),
    .A1(_1003_),
    .S(net10),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2086_ (.A0(net145),
    .A1(_1008_),
    .S(net10),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2087_ (.A0(net159),
    .A1(_1012_),
    .S(_0495_),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_4 _2088_ (.A(_0809_),
    .B(_0977_),
    .Y(_0496_));
 sky130_fd_sc_hd__mux2_1 _2089_ (.A0(net188),
    .A1(_0980_),
    .S(_0496_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2090_ (.A0(net171),
    .A1(_0987_),
    .S(_0496_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2091_ (.A0(net170),
    .A1(_0992_),
    .S(_0496_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2092_ (.A0(net148),
    .A1(_0996_),
    .S(_0496_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2093_ (.A0(net191),
    .A1(_0997_),
    .S(_0496_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(net158),
    .A1(_1003_),
    .S(_0496_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2095_ (.A0(net139),
    .A1(_1008_),
    .S(_0496_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(net184),
    .A1(_1012_),
    .S(_0496_),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _2097_ (.A1(net166),
    .A2(net33),
    .B1(net24),
    .B2(net168),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_1 _2098_ (.A1(\spi_sram_master_inst.data[25] ),
    .A2(net33),
    .B1(net23),
    .B2(net166),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _2099_ (.A1(net183),
    .A2(net33),
    .B1(net24),
    .B2(net187),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _2100_ (.A1(net169),
    .A2(net32),
    .B1(net23),
    .B2(net183),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _2101_ (.A1(net146),
    .A2(net32),
    .B1(net23),
    .B2(net169),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _2102_ (.A1(\spi_sram_master_inst.data[29] ),
    .A2(net32),
    .B1(net23),
    .B2(net146),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _2103_ (.A1(net133),
    .A2(net32),
    .B1(net23),
    .B2(net176),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _2104_ (.A1(\spi_sram_master_inst.data[31] ),
    .A2(net33),
    .B1(net24),
    .B2(net133),
    .X(_0170_));
 sky130_fd_sc_hd__o22a_1 _2105_ (.A1(net162),
    .A2(_0821_),
    .B1(_0823_),
    .B2(net165),
    .X(_0171_));
 sky130_fd_sc_hd__a22o_1 _2106_ (.A1(net155),
    .A2(net32),
    .B1(net23),
    .B2(net162),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_1 _2107_ (.A1(net151),
    .A2(net32),
    .B1(net23),
    .B2(net155),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_1 _2108_ (.A1(\spi_sram_master_inst.data[36] ),
    .A2(net32),
    .B1(net23),
    .B2(net151),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _2109_ (.A1(\spi_sram_master_inst.data[37] ),
    .A2(net32),
    .B1(net23),
    .B2(net156),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _2110_ (.A1(net131),
    .A2(net32),
    .B1(net23),
    .B2(net177),
    .X(_0176_));
 sky130_fd_sc_hd__o22a_1 _2111_ (.A1(\spi_sram_master_inst.data[39] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(net131),
    .X(_0177_));
 sky130_fd_sc_hd__o21ai_1 _2112_ (.A1(_1015_),
    .A2(_0278_),
    .B1(net63),
    .Y(_0497_));
 sky130_fd_sc_hd__o22a_1 _2113_ (.A1(net203),
    .A2(net63),
    .B1(_0280_),
    .B2(_0497_),
    .X(_0178_));
 sky130_fd_sc_hd__and3_4 _2114_ (.A(net16),
    .B(_0805_),
    .C(_0978_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(net163),
    .A1(_0980_),
    .S(_0498_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2116_ (.A0(net160),
    .A1(_0987_),
    .S(_0498_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(net174),
    .A1(_0992_),
    .S(_0498_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(net141),
    .A1(_0996_),
    .S(_0498_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2119_ (.A0(net192),
    .A1(_0997_),
    .S(_0498_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2120_ (.A0(net179),
    .A1(_1003_),
    .S(_0498_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2121_ (.A0(net182),
    .A1(_1008_),
    .S(_0498_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2122_ (.A0(net178),
    .A1(_1012_),
    .S(_0498_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _2124_ (.CLK(clknet_4_4_0_clk),
    .D(net128),
    .Q(\spi_sram_master_inst.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2125_ (.CLK(clknet_4_4_0_clk),
    .D(_0018_),
    .Q(\spi_sram_master_inst.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2126_ (.CLK(clknet_4_6_0_clk),
    .D(_0019_),
    .Q(\cpu_inst.DI[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2127_ (.CLK(clknet_4_12_0_clk),
    .D(_0020_),
    .Q(\cpu_inst.DI[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2128_ (.CLK(clknet_4_12_0_clk),
    .D(_0021_),
    .Q(\cpu_inst.DI[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2129_ (.CLK(clknet_4_9_0_clk),
    .D(_0022_),
    .Q(\cpu_inst.DI[3] ));
 sky130_fd_sc_hd__dfxtp_4 _2130_ (.CLK(clknet_4_12_0_clk),
    .D(_0023_),
    .Q(\cpu_inst.DI[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2131_ (.CLK(clknet_4_12_0_clk),
    .D(_0024_),
    .Q(\cpu_inst.DI[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2132_ (.CLK(clknet_4_9_0_clk),
    .D(_0025_),
    .Q(\cpu_inst.DI[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2133_ (.CLK(clknet_4_9_0_clk),
    .D(_0026_),
    .Q(\cpu_inst.DI[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2134_ (.CLK(clknet_4_15_0_clk),
    .D(_0027_),
    .Q(\spi_sram_master_inst.data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2135_ (.CLK(clknet_4_15_0_clk),
    .D(_0028_),
    .Q(\spi_sram_master_inst.data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2136_ (.CLK(clknet_4_15_0_clk),
    .D(_0029_),
    .Q(\spi_sram_master_inst.data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2137_ (.CLK(clknet_4_15_0_clk),
    .D(_0030_),
    .Q(\spi_sram_master_inst.data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2138_ (.CLK(clknet_4_15_0_clk),
    .D(_0031_),
    .Q(\spi_sram_master_inst.data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2139_ (.CLK(clknet_4_15_0_clk),
    .D(_0032_),
    .Q(\spi_sram_master_inst.data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2140_ (.CLK(clknet_4_15_0_clk),
    .D(_0033_),
    .Q(\spi_sram_master_inst.data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2141_ (.CLK(clknet_4_13_0_clk),
    .D(_0034_),
    .Q(\spi_sram_master_inst.data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2142_ (.CLK(clknet_4_13_0_clk),
    .D(_0035_),
    .Q(\spi_sram_master_inst.data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2143_ (.CLK(clknet_4_13_0_clk),
    .D(_0036_),
    .Q(\spi_sram_master_inst.data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2144_ (.CLK(clknet_4_13_0_clk),
    .D(_0037_),
    .Q(\spi_sram_master_inst.data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2145_ (.CLK(clknet_4_13_0_clk),
    .D(_0038_),
    .Q(\spi_sram_master_inst.data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2146_ (.CLK(clknet_4_13_0_clk),
    .D(_0039_),
    .Q(\spi_sram_master_inst.data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2147_ (.CLK(clknet_4_6_0_clk),
    .D(_0040_),
    .Q(\spi_sram_master_inst.data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2148_ (.CLK(clknet_4_6_0_clk),
    .D(_0041_),
    .Q(\spi_sram_master_inst.data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2149_ (.CLK(clknet_4_6_0_clk),
    .D(_0042_),
    .Q(\spi_sram_master_inst.data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2150_ (.CLK(clknet_4_6_0_clk),
    .D(_0043_),
    .Q(\spi_sram_master_inst.data[32] ));
 sky130_fd_sc_hd__dfrtp_1 _2151_ (.CLK(clknet_4_1_0_clk),
    .D(_0009_),
    .RESET_B(net101),
    .Q(\cpu_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2152_ (.CLK(clknet_4_1_0_clk),
    .D(_0010_),
    .RESET_B(net101),
    .Q(\cpu_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2153_ (.CLK(clknet_4_1_0_clk),
    .D(_0011_),
    .RESET_B(net101),
    .Q(\cpu_inst.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _2154_ (.CLK(clknet_4_1_0_clk),
    .D(_0012_),
    .SET_B(net101),
    .Q(\cpu_inst.state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2155_ (.CLK(clknet_4_1_0_clk),
    .D(_0013_),
    .RESET_B(net101),
    .Q(\cpu_inst.state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2156_ (.CLK(clknet_4_1_0_clk),
    .D(_0014_),
    .RESET_B(net101),
    .Q(\cpu_inst.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2157_ (.CLK(clknet_4_8_0_clk),
    .D(_0044_),
    .Q(\cpu_inst.AXYS[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2158_ (.CLK(clknet_4_10_0_clk),
    .D(_0045_),
    .Q(\cpu_inst.AXYS[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2159_ (.CLK(clknet_4_11_0_clk),
    .D(_0046_),
    .Q(\cpu_inst.AXYS[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2160_ (.CLK(clknet_4_10_0_clk),
    .D(_0047_),
    .Q(\cpu_inst.AXYS[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2161_ (.CLK(clknet_4_11_0_clk),
    .D(_0048_),
    .Q(\cpu_inst.AXYS[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2162_ (.CLK(clknet_4_8_0_clk),
    .D(_0049_),
    .Q(\cpu_inst.AXYS[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2163_ (.CLK(clknet_4_10_0_clk),
    .D(_0050_),
    .Q(\cpu_inst.AXYS[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2164_ (.CLK(clknet_4_8_0_clk),
    .D(_0051_),
    .Q(\cpu_inst.AXYS[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2165_ (.CLK(clknet_4_4_0_clk),
    .D(_0006_),
    .Q(\spi_sram_master_inst.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2166_ (.CLK(clknet_4_4_0_clk),
    .D(_0007_),
    .Q(\spi_sram_master_inst.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2167_ (.CLK(clknet_4_5_0_clk),
    .D(_0008_),
    .Q(\spi_sram_master_inst.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2168_ (.CLK(clknet_4_9_0_clk),
    .D(_0052_),
    .Q(\cpu_inst.backwards ));
 sky130_fd_sc_hd__dfxtp_1 _2169_ (.CLK(clknet_4_11_0_clk),
    .D(_0053_),
    .Q(\cpu_inst.ALU.CO ));
 sky130_fd_sc_hd__dfxtp_1 _2170_ (.CLK(clknet_4_14_0_clk),
    .D(_0054_),
    .Q(\cpu_inst.ADD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2171_ (.CLK(clknet_4_11_0_clk),
    .D(_0055_),
    .Q(\cpu_inst.ADD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2172_ (.CLK(clknet_4_11_0_clk),
    .D(_0056_),
    .Q(\cpu_inst.ADD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2173_ (.CLK(clknet_4_11_0_clk),
    .D(_0057_),
    .Q(\cpu_inst.ADD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2174_ (.CLK(clknet_4_11_0_clk),
    .D(_0058_),
    .Q(\cpu_inst.ADD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2175_ (.CLK(clknet_4_11_0_clk),
    .D(_0059_),
    .Q(\cpu_inst.ADD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2176_ (.CLK(clknet_4_11_0_clk),
    .D(_0060_),
    .Q(\cpu_inst.ADD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2177_ (.CLK(clknet_4_11_0_clk),
    .D(_0061_),
    .Q(\cpu_inst.ADD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2178_ (.CLK(clknet_4_11_0_clk),
    .D(_0062_),
    .Q(\cpu_inst.ALU.HC ));
 sky130_fd_sc_hd__dfxtp_1 _2179_ (.CLK(clknet_4_9_0_clk),
    .D(_0063_),
    .Q(\cpu_inst.ALU.AI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2180_ (.CLK(clknet_4_12_0_clk),
    .D(_0064_),
    .Q(\cpu_inst.ABH[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2181_ (.CLK(clknet_4_12_0_clk),
    .D(_0065_),
    .Q(\cpu_inst.ABH[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2182_ (.CLK(clknet_4_12_0_clk),
    .D(_0066_),
    .Q(\cpu_inst.ABH[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2183_ (.CLK(clknet_4_13_0_clk),
    .D(_0067_),
    .Q(\cpu_inst.ABH[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2184_ (.CLK(clknet_4_13_0_clk),
    .D(_0068_),
    .Q(\cpu_inst.ABH[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2185_ (.CLK(clknet_4_13_0_clk),
    .D(_0069_),
    .Q(\cpu_inst.ABH[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2186_ (.CLK(clknet_4_6_0_clk),
    .D(_0070_),
    .Q(\cpu_inst.ABH[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2187_ (.CLK(clknet_4_6_0_clk),
    .D(_0071_),
    .Q(\cpu_inst.ABH[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2188_ (.CLK(clknet_4_14_0_clk),
    .D(_0072_),
    .Q(\cpu_inst.ABL[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2189_ (.CLK(clknet_4_14_0_clk),
    .D(_0073_),
    .Q(\cpu_inst.ABL[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2190_ (.CLK(clknet_4_14_0_clk),
    .D(_0074_),
    .Q(\cpu_inst.ABL[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2191_ (.CLK(clknet_4_15_0_clk),
    .D(_0075_),
    .Q(\cpu_inst.ABL[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2192_ (.CLK(clknet_4_15_0_clk),
    .D(_0076_),
    .Q(\cpu_inst.ABL[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2193_ (.CLK(clknet_4_15_0_clk),
    .D(_0077_),
    .Q(\cpu_inst.ABL[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2194_ (.CLK(clknet_4_14_0_clk),
    .D(_0078_),
    .Q(\cpu_inst.ABL[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2195_ (.CLK(clknet_4_13_0_clk),
    .D(_0079_),
    .Q(\cpu_inst.ABL[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2196_ (.CLK(clknet_4_9_0_clk),
    .D(_0080_),
    .Q(\cpu_inst.adj_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2197_ (.CLK(clknet_4_3_0_clk),
    .D(_0081_),
    .Q(\cpu_inst.C ));
 sky130_fd_sc_hd__dfxtp_1 _2198_ (.CLK(clknet_4_9_0_clk),
    .D(_0082_),
    .Q(\cpu_inst.Z ));
 sky130_fd_sc_hd__dfxtp_1 _2199_ (.CLK(clknet_4_9_0_clk),
    .D(_0083_),
    .Q(\cpu_inst.N ));
 sky130_fd_sc_hd__dfxtp_1 _2200_ (.CLK(clknet_4_9_0_clk),
    .D(_0084_),
    .Q(\cpu_inst.D ));
 sky130_fd_sc_hd__dfxtp_1 _2201_ (.CLK(clknet_4_3_0_clk),
    .D(_0085_),
    .Q(\cpu_inst.I ));
 sky130_fd_sc_hd__dfxtp_1 _2202_ (.CLK(clknet_4_9_0_clk),
    .D(_0086_),
    .Q(\cpu_inst.V ));
 sky130_fd_sc_hd__dfrtp_1 _2203_ (.CLK(clknet_4_8_0_clk),
    .D(_0087_),
    .RESET_B(net102),
    .Q(\cpu_inst.IRHOLD_valid ));
 sky130_fd_sc_hd__dfxtp_1 _2204_ (.CLK(clknet_4_8_0_clk),
    .D(_0088_),
    .Q(\cpu_inst.IRHOLD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2205_ (.CLK(clknet_4_8_0_clk),
    .D(_0089_),
    .Q(\cpu_inst.IRHOLD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2206_ (.CLK(clknet_4_8_0_clk),
    .D(_0090_),
    .Q(\cpu_inst.IRHOLD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2207_ (.CLK(clknet_4_9_0_clk),
    .D(_0091_),
    .Q(\cpu_inst.IRHOLD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2208_ (.CLK(clknet_4_8_0_clk),
    .D(_0092_),
    .Q(\cpu_inst.IRHOLD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2209_ (.CLK(clknet_4_8_0_clk),
    .D(_0093_),
    .Q(\cpu_inst.IRHOLD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2210_ (.CLK(clknet_4_8_0_clk),
    .D(_0094_),
    .Q(\cpu_inst.IRHOLD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2211_ (.CLK(clknet_4_8_0_clk),
    .D(_0095_),
    .Q(\cpu_inst.IRHOLD[7] ));
 sky130_fd_sc_hd__dfstp_1 _2212_ (.CLK(clknet_4_6_0_clk),
    .D(_0096_),
    .SET_B(net102),
    .Q(\cpu_inst.res ));
 sky130_fd_sc_hd__dfxtp_1 _2213_ (.CLK(clknet_4_0_0_clk),
    .D(_0097_),
    .Q(\cpu_inst.load_reg ));
 sky130_fd_sc_hd__dfxtp_1 _2214_ (.CLK(clknet_4_1_0_clk),
    .D(_0098_),
    .Q(\cpu_inst.dst_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2215_ (.CLK(clknet_4_2_0_clk),
    .D(_0099_),
    .Q(\cpu_inst.dst_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2216_ (.CLK(clknet_4_2_0_clk),
    .D(_0100_),
    .Q(\cpu_inst.src_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2217_ (.CLK(clknet_4_2_0_clk),
    .D(_0101_),
    .Q(\cpu_inst.src_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2218_ (.CLK(clknet_4_0_0_clk),
    .D(_0102_),
    .Q(\cpu_inst.index_y ));
 sky130_fd_sc_hd__dfxtp_1 _2219_ (.CLK(clknet_4_0_0_clk),
    .D(_0103_),
    .Q(\cpu_inst.store ));
 sky130_fd_sc_hd__dfxtp_1 _2220_ (.CLK(clknet_4_0_0_clk),
    .D(_0104_),
    .Q(\cpu_inst.write_back ));
 sky130_fd_sc_hd__dfxtp_1 _2221_ (.CLK(clknet_4_2_0_clk),
    .D(_0105_),
    .Q(\cpu_inst.load_only ));
 sky130_fd_sc_hd__dfxtp_1 _2222_ (.CLK(clknet_4_0_0_clk),
    .D(_0106_),
    .Q(\cpu_inst.inc ));
 sky130_fd_sc_hd__dfxtp_1 _2223_ (.CLK(clknet_4_3_0_clk),
    .D(_0107_),
    .Q(\cpu_inst.adc_sbc ));
 sky130_fd_sc_hd__dfxtp_1 _2224_ (.CLK(clknet_4_3_0_clk),
    .D(_0108_),
    .Q(\cpu_inst.shift ));
 sky130_fd_sc_hd__dfxtp_1 _2225_ (.CLK(clknet_4_3_0_clk),
    .D(_0109_),
    .Q(\cpu_inst.adc_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2226_ (.CLK(clknet_4_2_0_clk),
    .D(_0110_),
    .Q(\cpu_inst.compare ));
 sky130_fd_sc_hd__dfxtp_1 _2227_ (.CLK(clknet_4_3_0_clk),
    .D(_0111_),
    .Q(\cpu_inst.shift_right ));
 sky130_fd_sc_hd__dfxtp_1 _2228_ (.CLK(clknet_4_3_0_clk),
    .D(_0112_),
    .Q(\cpu_inst.rotate ));
 sky130_fd_sc_hd__dfxtp_1 _2229_ (.CLK(clknet_4_2_0_clk),
    .D(_0113_),
    .Q(\cpu_inst.op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2230_ (.CLK(clknet_4_3_0_clk),
    .D(_0114_),
    .Q(\cpu_inst.op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2231_ (.CLK(clknet_4_9_0_clk),
    .D(_0115_),
    .Q(\cpu_inst.op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2232_ (.CLK(clknet_4_2_0_clk),
    .D(_0116_),
    .Q(\cpu_inst.op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2233_ (.CLK(clknet_4_8_0_clk),
    .D(_0117_),
    .Q(\cpu_inst.bit_ins ));
 sky130_fd_sc_hd__dfxtp_1 _2234_ (.CLK(clknet_4_2_0_clk),
    .D(_0118_),
    .Q(\cpu_inst.clv ));
 sky130_fd_sc_hd__dfxtp_1 _2235_ (.CLK(clknet_4_2_0_clk),
    .D(_0119_),
    .Q(\cpu_inst.sei ));
 sky130_fd_sc_hd__dfxtp_1 _2236_ (.CLK(clknet_4_2_0_clk),
    .D(_0120_),
    .Q(\cpu_inst.cli ));
 sky130_fd_sc_hd__dfxtp_1 _2237_ (.CLK(clknet_4_2_0_clk),
    .D(_0121_),
    .Q(\cpu_inst.sed ));
 sky130_fd_sc_hd__dfxtp_1 _2238_ (.CLK(clknet_4_8_0_clk),
    .D(_0122_),
    .Q(\cpu_inst.cld ));
 sky130_fd_sc_hd__dfxtp_1 _2239_ (.CLK(clknet_4_2_0_clk),
    .D(_0123_),
    .Q(\cpu_inst.sec ));
 sky130_fd_sc_hd__dfxtp_1 _2240_ (.CLK(clknet_4_2_0_clk),
    .D(_0124_),
    .Q(\cpu_inst.clc ));
 sky130_fd_sc_hd__dfxtp_1 _2241_ (.CLK(clknet_4_0_0_clk),
    .D(_0125_),
    .Q(\cpu_inst.php ));
 sky130_fd_sc_hd__dfxtp_1 _2242_ (.CLK(clknet_4_0_0_clk),
    .D(_0126_),
    .Q(\cpu_inst.plp ));
 sky130_fd_sc_hd__dfxtp_1 _2243_ (.CLK(clknet_4_1_0_clk),
    .D(_0127_),
    .Q(\cpu_inst.cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2244_ (.CLK(clknet_4_9_0_clk),
    .D(_0128_),
    .Q(\cpu_inst.cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2245_ (.CLK(clknet_4_8_0_clk),
    .D(_0129_),
    .Q(\cpu_inst.cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2246_ (.CLK(clknet_4_14_0_clk),
    .D(_0130_),
    .Q(\cpu_inst.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2247_ (.CLK(clknet_4_14_0_clk),
    .D(_0131_),
    .Q(\cpu_inst.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2248_ (.CLK(clknet_4_14_0_clk),
    .D(_0132_),
    .Q(\cpu_inst.PC[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2249_ (.CLK(clknet_4_15_0_clk),
    .D(_0133_),
    .Q(\cpu_inst.PC[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2250_ (.CLK(clknet_4_15_0_clk),
    .D(_0134_),
    .Q(\cpu_inst.PC[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2251_ (.CLK(clknet_4_14_0_clk),
    .D(_0135_),
    .Q(\cpu_inst.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2252_ (.CLK(clknet_4_14_0_clk),
    .D(_0136_),
    .Q(\cpu_inst.PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2253_ (.CLK(clknet_4_12_0_clk),
    .D(_0137_),
    .Q(\cpu_inst.PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2254_ (.CLK(clknet_4_13_0_clk),
    .D(_0138_),
    .Q(\cpu_inst.PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2255_ (.CLK(clknet_4_13_0_clk),
    .D(_0139_),
    .Q(\cpu_inst.PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2256_ (.CLK(clknet_4_12_0_clk),
    .D(_0140_),
    .Q(\cpu_inst.PC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2257_ (.CLK(clknet_4_12_0_clk),
    .D(_0141_),
    .Q(\cpu_inst.PC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2258_ (.CLK(clknet_4_13_0_clk),
    .D(_0142_),
    .Q(\cpu_inst.PC[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2259_ (.CLK(clknet_4_6_0_clk),
    .D(_0143_),
    .Q(\cpu_inst.PC[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2260_ (.CLK(clknet_4_6_0_clk),
    .D(_0144_),
    .Q(\cpu_inst.PC[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2261_ (.CLK(clknet_4_6_0_clk),
    .D(_0145_),
    .Q(\cpu_inst.PC[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2262_ (.CLK(clknet_4_7_0_clk),
    .D(net3),
    .Q(\cpu_inst.NMI_1 ));
 sky130_fd_sc_hd__dfxtp_1 _2263_ (.CLK(clknet_4_7_0_clk),
    .D(_0146_),
    .Q(\cpu_inst.NMI_edge ));
 sky130_fd_sc_hd__dfstp_1 _2264_ (.CLK(clknet_4_5_0_clk),
    .D(net103),
    .SET_B(net101),
    .Q(\spi_sram_master_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2265_ (.CLK(clknet_4_4_0_clk),
    .D(_0000_),
    .RESET_B(net101),
    .Q(\spi_sram_master_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2266_ (.CLK(clknet_4_4_0_clk),
    .D(_0001_),
    .RESET_B(net101),
    .Q(\spi_sram_master_inst.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2267_ (.CLK(clknet_4_5_0_clk),
    .D(_0002_),
    .RESET_B(net101),
    .Q(\spi_sram_master_inst.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2268_ (.CLK(clknet_4_4_0_clk),
    .D(_0004_),
    .RESET_B(net102),
    .Q(\spi_sram_master_inst.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2269_ (.CLK(clknet_4_5_0_clk),
    .D(net129),
    .RESET_B(net102),
    .Q(\spi_sram_master_inst.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2270_ (.CLK(clknet_4_4_0_clk),
    .D(net210),
    .RESET_B(net102),
    .Q(\spi_sram_master_inst.state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2271_ (.CLK(clknet_4_5_0_clk),
    .D(net208),
    .RESET_B(net102),
    .Q(\spi_sram_master_inst.state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2272_ (.CLK(clknet_4_8_0_clk),
    .D(_0147_),
    .Q(\cpu_inst.AXYS[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2273_ (.CLK(clknet_4_10_0_clk),
    .D(_0148_),
    .Q(\cpu_inst.AXYS[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2274_ (.CLK(clknet_4_10_0_clk),
    .D(_0149_),
    .Q(\cpu_inst.AXYS[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2275_ (.CLK(clknet_4_10_0_clk),
    .D(_0150_),
    .Q(\cpu_inst.AXYS[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2276_ (.CLK(clknet_4_10_0_clk),
    .D(_0151_),
    .Q(\cpu_inst.AXYS[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2277_ (.CLK(clknet_4_8_0_clk),
    .D(_0152_),
    .Q(\cpu_inst.AXYS[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2278_ (.CLK(clknet_4_10_0_clk),
    .D(_0153_),
    .Q(\cpu_inst.AXYS[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2279_ (.CLK(clknet_4_8_0_clk),
    .D(_0154_),
    .Q(\cpu_inst.AXYS[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2280_ (.CLK(clknet_4_8_0_clk),
    .D(_0155_),
    .Q(\cpu_inst.AXYS[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2281_ (.CLK(clknet_4_10_0_clk),
    .D(_0156_),
    .Q(\cpu_inst.AXYS[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2282_ (.CLK(clknet_4_11_0_clk),
    .D(_0157_),
    .Q(\cpu_inst.AXYS[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2283_ (.CLK(clknet_4_10_0_clk),
    .D(_0158_),
    .Q(\cpu_inst.AXYS[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2284_ (.CLK(clknet_4_11_0_clk),
    .D(_0159_),
    .Q(\cpu_inst.AXYS[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2285_ (.CLK(clknet_4_8_0_clk),
    .D(_0160_),
    .Q(\cpu_inst.AXYS[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2286_ (.CLK(clknet_4_10_0_clk),
    .D(_0161_),
    .Q(\cpu_inst.AXYS[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2287_ (.CLK(clknet_4_8_0_clk),
    .D(_0162_),
    .Q(\cpu_inst.AXYS[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2288_ (.CLK(clknet_4_6_0_clk),
    .D(_0163_),
    .Q(\spi_sram_master_inst.data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2289_ (.CLK(clknet_4_6_0_clk),
    .D(net167),
    .Q(\spi_sram_master_inst.data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2290_ (.CLK(clknet_4_7_0_clk),
    .D(_0165_),
    .Q(\spi_sram_master_inst.data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2291_ (.CLK(clknet_4_7_0_clk),
    .D(_0166_),
    .Q(\spi_sram_master_inst.data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2292_ (.CLK(clknet_4_7_0_clk),
    .D(_0167_),
    .Q(\spi_sram_master_inst.data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2293_ (.CLK(clknet_4_7_0_clk),
    .D(net147),
    .Q(\spi_sram_master_inst.data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2294_ (.CLK(clknet_4_7_0_clk),
    .D(_0169_),
    .Q(\spi_sram_master_inst.data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2295_ (.CLK(clknet_4_6_0_clk),
    .D(net134),
    .Q(\spi_sram_master_inst.data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2296_ (.CLK(clknet_4_5_0_clk),
    .D(_0171_),
    .Q(\spi_sram_master_inst.data[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2297_ (.CLK(clknet_4_7_0_clk),
    .D(_0172_),
    .Q(\spi_sram_master_inst.data[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2298_ (.CLK(clknet_4_7_0_clk),
    .D(_0173_),
    .Q(\spi_sram_master_inst.data[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2299_ (.CLK(clknet_4_7_0_clk),
    .D(net152),
    .Q(\spi_sram_master_inst.data[36] ));
 sky130_fd_sc_hd__dfxtp_1 _2300_ (.CLK(clknet_4_7_0_clk),
    .D(net157),
    .Q(\spi_sram_master_inst.data[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2301_ (.CLK(clknet_4_7_0_clk),
    .D(_0176_),
    .Q(\spi_sram_master_inst.data[38] ));
 sky130_fd_sc_hd__dfxtp_1 _2302_ (.CLK(clknet_4_7_0_clk),
    .D(net132),
    .Q(\spi_sram_master_inst.data[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2303_ (.CLK(clknet_4_9_0_clk),
    .D(_0178_),
    .Q(\cpu_inst.ALU.BI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2304_ (.CLK(net125),
    .D(\spi_sram_master_inst.data[39] ),
    .Q(\spi_sram_master_inst.dout ));
 sky130_fd_sc_hd__dfxtp_1 _2305_ (.CLK(net126),
    .D(\spi_sram_master_inst.cs_n_sm ),
    .Q(\spi_sram_master_inst.cs_n ));
 sky130_fd_sc_hd__dfxtp_1 _2306_ (.CLK(clknet_4_8_0_clk),
    .D(_0179_),
    .Q(\cpu_inst.AXYS[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2307_ (.CLK(clknet_4_10_0_clk),
    .D(_0180_),
    .Q(\cpu_inst.AXYS[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2308_ (.CLK(clknet_4_11_0_clk),
    .D(_0181_),
    .Q(\cpu_inst.AXYS[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2309_ (.CLK(clknet_4_10_0_clk),
    .D(_0182_),
    .Q(\cpu_inst.AXYS[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2310_ (.CLK(clknet_4_10_0_clk),
    .D(_0183_),
    .Q(\cpu_inst.AXYS[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2311_ (.CLK(clknet_4_8_0_clk),
    .D(_0184_),
    .Q(\cpu_inst.AXYS[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2312_ (.CLK(clknet_4_10_0_clk),
    .D(_0185_),
    .Q(\cpu_inst.AXYS[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2313_ (.CLK(clknet_4_8_0_clk),
    .D(_0186_),
    .Q(\cpu_inst.AXYS[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2314_ (.CLK(clknet_4_5_0_clk),
    .D(_0187_),
    .Q(\spi_sram_master_inst.counter_done ));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_124 (.HI(net124));
 sky130_fd_sc_hd__inv_2 _1074__1 (.A(clknet_4_5_0_clk),
    .Y(net125));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_122 (.HI(net122));
 sky130_fd_sc_hd__buf_2 _2337_ (.A(\spi_sram_master_inst.cs_n ),
    .X(uio_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _2338_ (.A(\spi_sram_master_inst.dout ),
    .X(uio_out[1]));
 sky130_fd_sc_hd__buf_2 _2339_ (.A(clknet_4_5_0_clk),
    .X(uio_out[3]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1198 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[6]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[7]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(uio_in[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 fanout5 (.A(_0304_),
    .X(net5));
 sky130_fd_sc_hd__buf_2 fanout6 (.A(_0304_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net9),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 fanout8 (.A(_0897_),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 max_cap9 (.A(_0897_),
    .X(net9));
 sky130_fd_sc_hd__buf_2 max_cap10 (.A(_0495_),
    .X(net10));
 sky130_fd_sc_hd__buf_1 wire11 (.A(_0396_),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 max_cap12 (.A(_1024_),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(_1014_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 max_cap15 (.A(_0805_),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(_0803_),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(_0803_),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(_0298_),
    .X(net19));
 sky130_fd_sc_hd__buf_1 max_cap20 (.A(_0796_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(_0414_),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(_0414_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(_0822_),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(_0822_),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(_0542_),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(_0541_),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_1 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout34 (.A(net36),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(_0820_),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(_0670_),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(_0632_),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net41),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(_0582_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(_0578_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(_0571_),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(_0566_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(_0540_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(_0539_),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(_0530_),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(_0560_),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(_0560_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(_0536_),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(_0525_),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(_0525_),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net58),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net67),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net67),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(net67),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net66),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(_0523_),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net71),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(_0522_),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(_0522_),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(\cpu_inst.plp ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(\cpu_inst.IRHOLD_valid ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(\cpu_inst.ADD[7] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(\cpu_inst.ADD[6] ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(\cpu_inst.ADD[5] ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(\cpu_inst.ADD[4] ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(\cpu_inst.ADD[3] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(\cpu_inst.ADD[2] ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(\cpu_inst.ADD[1] ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(\cpu_inst.ADD[0] ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(\cpu_inst.ALU.CO ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(\cpu_inst.state[5] ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(\cpu_inst.state[4] ),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(\cpu_inst.state[3] ),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(\cpu_inst.state[2] ),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(\cpu_inst.state[2] ),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(\cpu_inst.state[1] ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(\cpu_inst.state[1] ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 fanout93 (.A(\cpu_inst.state[0] ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(\cpu_inst.state[0] ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(\cpu_inst.DI[7] ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(\cpu_inst.DI[6] ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 fanout97 (.A(\cpu_inst.DI[3] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(\cpu_inst.DI[2] ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(\cpu_inst.DI[1] ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 fanout100 (.A(\cpu_inst.DI[0] ),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(net1),
    .X(net102));
 sky130_fd_sc_hd__conb_1 _2264__103 (.LO(net103));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__inv_12 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_12 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__inv_8 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_12 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__inv_12 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__inv_8 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__inv_8 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_8 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__inv_8 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__inv_8 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_12 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_8 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__inv_12 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\spi_sram_master_inst.counter[0] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0017_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\spi_sram_master_inst.state[1] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\spi_sram_master_inst.counter[4] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\spi_sram_master_inst.data[38] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0177_),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\spi_sram_master_inst.data[30] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0170_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\cpu_inst.AXYS[3][4] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\cpu_inst.dst_reg[1] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\cpu_inst.AXYS[3][3] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\cpu_inst.sec ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\cpu_inst.AXYS[1][6] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\cpu_inst.IRHOLD[1] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\cpu_inst.AXYS[0][3] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\cpu_inst.AXYS[3][5] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\cpu_inst.AXYS[3][2] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\cpu_inst.AXYS[3][1] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\cpu_inst.AXYS[3][6] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\spi_sram_master_inst.data[28] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0168_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\cpu_inst.AXYS[1][3] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\cpu_inst.IRHOLD[3] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\cpu_inst.op[2] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\spi_sram_master_inst.data[35] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0174_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\cpu_inst.IRHOLD[6] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\cpu_inst.IRHOLD[0] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\spi_sram_master_inst.data[34] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\spi_sram_master_inst.data[36] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0175_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\cpu_inst.AXYS[1][5] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\cpu_inst.AXYS[3][7] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\cpu_inst.AXYS[0][1] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\cpu_inst.IRHOLD[4] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\spi_sram_master_inst.data[33] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\cpu_inst.AXYS[0][0] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\cpu_inst.IRHOLD[7] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\spi_sram_master_inst.data[32] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\spi_sram_master_inst.data[24] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0164_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\spi_sram_master_inst.data[23] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\spi_sram_master_inst.data[27] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\cpu_inst.AXYS[1][2] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\cpu_inst.AXYS[1][1] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\cpu_inst.AXYS[2][3] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\cpu_inst.IRHOLD[2] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\cpu_inst.AXYS[0][2] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\cpu_inst.DI[1] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\spi_sram_master_inst.data[29] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\spi_sram_master_inst.data[37] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\cpu_inst.AXYS[0][7] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\cpu_inst.AXYS[0][5] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\cpu_inst.AXYS[2][7] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\cpu_inst.AXYS[2][5] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\cpu_inst.AXYS[0][6] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\spi_sram_master_inst.data[26] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\cpu_inst.AXYS[1][7] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\cpu_inst.AXYS[2][2] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\cpu_inst.AXYS[2][1] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\spi_sram_master_inst.data[25] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\cpu_inst.AXYS[1][0] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\cpu_inst.AXYS[2][6] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\cpu_inst.sed ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\cpu_inst.AXYS[1][4] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\cpu_inst.AXYS[0][4] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\cpu_inst.AXYS[2][4] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\cpu_inst.ADD[0] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\cpu_inst.index_y ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\cpu_inst.src_reg[0] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\cpu_inst.ALU.AI7 ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\cpu_inst.inc ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\cpu_inst.AXYS[3][0] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\cpu_inst.cond_code[2] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\spi_sram_master_inst.counter[1] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\cpu_inst.cond_code[0] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\cpu_inst.ALU.BI7 ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\cpu_inst.ABL[5] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\cpu_inst.NMI_1 ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\cpu_inst.ABL[6] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\spi_sram_master_inst.counter_done ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0003_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\spi_sram_master_inst.state[6] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0005_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\cpu_inst.PC[13] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\cpu_inst.ALU.HC ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\cpu_inst.ABL[1] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\cpu_inst.ABL[0] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\spi_sram_master_inst.data[31] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\cpu_inst.ABL[7] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\cpu_inst.V ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\cpu_inst.ABL[2] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\cpu_inst.AXYS[2][0] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\cpu_inst.ABL[4] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\spi_sram_master_inst.state[3] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\cpu_inst.N ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\spi_sram_master_inst.state[4] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\cpu_inst.PC[8] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\cpu_inst.cond_code[1] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\spi_sram_master_inst.counter_done ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\cpu_inst.ABL[3] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\cpu_inst.rotate ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\cpu_inst.ABH[6] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\cpu_inst.ABH[0] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\cpu_inst.clc ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\spi_sram_master_inst.state[7] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\cpu_inst.ABH[3] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\cpu_inst.ABH[2] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\cpu_inst.ABH[7] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\cpu_inst.ABH[5] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\cpu_inst.IRHOLD[5] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\cpu_inst.Z ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\cpu_inst.cli ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\cpu_inst.ABH[4] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\cpu_inst.PC[4] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\cpu_inst.adj_bcd ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\cpu_inst.load_only ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\cpu_inst.shift ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\cpu_inst.res ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\cpu_inst.ABH[1] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\cpu_inst.clv ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\cpu_inst.load_reg ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\spi_sram_master_inst.data[17] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\cpu_inst.bit_ins ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\spi_sram_master_inst.data[12] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0928_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\cpu_inst.PC[11] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\cpu_inst.I ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\spi_sram_master_inst.data[8] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0908_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\cpu_inst.compare ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\spi_sram_master_inst.data[20] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0964_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\spi_sram_master_inst.data[20] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0960_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\spi_sram_master_inst.data[9] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\spi_sram_master_inst.data[13] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0933_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\spi_sram_master_inst.data[10] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\spi_sram_master_inst.data[21] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0968_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\spi_sram_master_inst.data[14] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\cpu_inst.PC[15] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\cpu_inst.PC[10] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\spi_sram_master_inst.data[22] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\spi_sram_master_inst.data[19] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0956_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\cpu_inst.PC[9] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\spi_sram_master_inst.data[16] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0944_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\cpu_inst.cld ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\spi_sram_master_inst.data[11] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\cpu_inst.PC[12] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\spi_sram_master_inst.data[10] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\spi_sram_master_inst.data[16] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0948_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\spi_sram_master_inst.data[11] ),
    .X(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net46));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 assign uio_oe[0] = net122;
 assign uio_oe[1] = net123;
 assign uio_oe[2] = net104;
 assign uio_oe[3] = net124;
 assign uio_oe[4] = net105;
 assign uio_oe[5] = net106;
 assign uio_oe[6] = net107;
 assign uio_oe[7] = net108;
 assign uio_out[2] = net109;
 assign uio_out[4] = net110;
 assign uio_out[5] = net111;
 assign uio_out[6] = net112;
 assign uio_out[7] = net113;
 assign uo_out[0] = net114;
 assign uo_out[1] = net115;
 assign uo_out[2] = net116;
 assign uo_out[3] = net117;
 assign uo_out[4] = net118;
 assign uo_out[5] = net119;
 assign uo_out[6] = net120;
 assign uo_out[7] = net121;
endmodule
