module tt_um_anders_tt_6502 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire net123;
 wire clknet_0_clk;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire \cpu_inst.ABH[0] ;
 wire \cpu_inst.ABH[1] ;
 wire \cpu_inst.ABH[2] ;
 wire \cpu_inst.ABH[3] ;
 wire \cpu_inst.ABH[4] ;
 wire \cpu_inst.ABH[5] ;
 wire \cpu_inst.ABH[6] ;
 wire \cpu_inst.ABH[7] ;
 wire \cpu_inst.ABL[0] ;
 wire \cpu_inst.ABL[1] ;
 wire \cpu_inst.ABL[2] ;
 wire \cpu_inst.ABL[3] ;
 wire \cpu_inst.ABL[4] ;
 wire \cpu_inst.ABL[5] ;
 wire \cpu_inst.ABL[6] ;
 wire \cpu_inst.ABL[7] ;
 wire \cpu_inst.ADD[0] ;
 wire \cpu_inst.ADD[1] ;
 wire \cpu_inst.ADD[2] ;
 wire \cpu_inst.ADD[3] ;
 wire \cpu_inst.ADD[4] ;
 wire \cpu_inst.ADD[5] ;
 wire \cpu_inst.ADD[6] ;
 wire \cpu_inst.ADD[7] ;
 wire \cpu_inst.ALU.AI7 ;
 wire \cpu_inst.ALU.BI7 ;
 wire \cpu_inst.ALU.CO ;
 wire \cpu_inst.ALU.HC ;
 wire \cpu_inst.AXYS[0][0] ;
 wire \cpu_inst.AXYS[0][1] ;
 wire \cpu_inst.AXYS[0][2] ;
 wire \cpu_inst.AXYS[0][3] ;
 wire \cpu_inst.AXYS[0][4] ;
 wire \cpu_inst.AXYS[0][5] ;
 wire \cpu_inst.AXYS[0][6] ;
 wire \cpu_inst.AXYS[0][7] ;
 wire \cpu_inst.AXYS[1][0] ;
 wire \cpu_inst.AXYS[1][1] ;
 wire \cpu_inst.AXYS[1][2] ;
 wire \cpu_inst.AXYS[1][3] ;
 wire \cpu_inst.AXYS[1][4] ;
 wire \cpu_inst.AXYS[1][5] ;
 wire \cpu_inst.AXYS[1][6] ;
 wire \cpu_inst.AXYS[1][7] ;
 wire \cpu_inst.AXYS[2][0] ;
 wire \cpu_inst.AXYS[2][1] ;
 wire \cpu_inst.AXYS[2][2] ;
 wire \cpu_inst.AXYS[2][3] ;
 wire \cpu_inst.AXYS[2][4] ;
 wire \cpu_inst.AXYS[2][5] ;
 wire \cpu_inst.AXYS[2][6] ;
 wire \cpu_inst.AXYS[2][7] ;
 wire \cpu_inst.AXYS[3][0] ;
 wire \cpu_inst.AXYS[3][1] ;
 wire \cpu_inst.AXYS[3][2] ;
 wire \cpu_inst.AXYS[3][3] ;
 wire \cpu_inst.AXYS[3][4] ;
 wire \cpu_inst.AXYS[3][5] ;
 wire \cpu_inst.AXYS[3][6] ;
 wire \cpu_inst.AXYS[3][7] ;
 wire \cpu_inst.C ;
 wire \cpu_inst.D ;
 wire \cpu_inst.DI[0] ;
 wire \cpu_inst.DI[1] ;
 wire \cpu_inst.DI[2] ;
 wire \cpu_inst.DI[3] ;
 wire \cpu_inst.DI[4] ;
 wire \cpu_inst.DI[5] ;
 wire \cpu_inst.DI[6] ;
 wire \cpu_inst.DI[7] ;
 wire \cpu_inst.I ;
 wire \cpu_inst.IRHOLD[0] ;
 wire \cpu_inst.IRHOLD[1] ;
 wire \cpu_inst.IRHOLD[2] ;
 wire \cpu_inst.IRHOLD[3] ;
 wire \cpu_inst.IRHOLD[4] ;
 wire \cpu_inst.IRHOLD[5] ;
 wire \cpu_inst.IRHOLD[6] ;
 wire \cpu_inst.IRHOLD[7] ;
 wire \cpu_inst.IRHOLD_valid ;
 wire \cpu_inst.N ;
 wire \cpu_inst.NMI_1 ;
 wire \cpu_inst.NMI_edge ;
 wire \cpu_inst.PC[0] ;
 wire \cpu_inst.PC[10] ;
 wire \cpu_inst.PC[11] ;
 wire \cpu_inst.PC[12] ;
 wire \cpu_inst.PC[13] ;
 wire \cpu_inst.PC[14] ;
 wire \cpu_inst.PC[15] ;
 wire \cpu_inst.PC[1] ;
 wire \cpu_inst.PC[2] ;
 wire \cpu_inst.PC[3] ;
 wire \cpu_inst.PC[4] ;
 wire \cpu_inst.PC[5] ;
 wire \cpu_inst.PC[6] ;
 wire \cpu_inst.PC[7] ;
 wire \cpu_inst.PC[8] ;
 wire \cpu_inst.PC[9] ;
 wire \cpu_inst.V ;
 wire \cpu_inst.Z ;
 wire \cpu_inst.adc_bcd ;
 wire \cpu_inst.adc_sbc ;
 wire \cpu_inst.adj_bcd ;
 wire \cpu_inst.backwards ;
 wire \cpu_inst.bit_ins ;
 wire \cpu_inst.clc ;
 wire \cpu_inst.cld ;
 wire \cpu_inst.cli ;
 wire \cpu_inst.clv ;
 wire \cpu_inst.compare ;
 wire \cpu_inst.cond_code[0] ;
 wire \cpu_inst.cond_code[1] ;
 wire \cpu_inst.cond_code[2] ;
 wire \cpu_inst.dst_reg[0] ;
 wire \cpu_inst.dst_reg[1] ;
 wire \cpu_inst.inc ;
 wire \cpu_inst.index_y ;
 wire \cpu_inst.load_only ;
 wire \cpu_inst.load_reg ;
 wire \cpu_inst.op[0] ;
 wire \cpu_inst.op[1] ;
 wire \cpu_inst.op[2] ;
 wire \cpu_inst.op[3] ;
 wire \cpu_inst.php ;
 wire \cpu_inst.plp ;
 wire \cpu_inst.res ;
 wire \cpu_inst.rotate ;
 wire \cpu_inst.sec ;
 wire \cpu_inst.sed ;
 wire \cpu_inst.sei ;
 wire \cpu_inst.shift ;
 wire \cpu_inst.shift_right ;
 wire \cpu_inst.src_reg[0] ;
 wire \cpu_inst.src_reg[1] ;
 wire \cpu_inst.state[0] ;
 wire \cpu_inst.state[1] ;
 wire \cpu_inst.state[2] ;
 wire \cpu_inst.state[3] ;
 wire \cpu_inst.state[4] ;
 wire \cpu_inst.state[5] ;
 wire \cpu_inst.store ;
 wire \cpu_inst.write_back ;
 wire \spi_sram_master_inst.counter[0] ;
 wire \spi_sram_master_inst.counter[1] ;
 wire \spi_sram_master_inst.counter[2] ;
 wire \spi_sram_master_inst.counter[3] ;
 wire \spi_sram_master_inst.counter[4] ;
 wire \spi_sram_master_inst.counter_done ;
 wire \spi_sram_master_inst.cs_n ;
 wire \spi_sram_master_inst.cs_n_sm ;
 wire \spi_sram_master_inst.data[10] ;
 wire \spi_sram_master_inst.data[11] ;
 wire \spi_sram_master_inst.data[12] ;
 wire \spi_sram_master_inst.data[13] ;
 wire \spi_sram_master_inst.data[14] ;
 wire \spi_sram_master_inst.data[15] ;
 wire \spi_sram_master_inst.data[16] ;
 wire \spi_sram_master_inst.data[17] ;
 wire \spi_sram_master_inst.data[18] ;
 wire \spi_sram_master_inst.data[19] ;
 wire \spi_sram_master_inst.data[20] ;
 wire \spi_sram_master_inst.data[21] ;
 wire \spi_sram_master_inst.data[22] ;
 wire \spi_sram_master_inst.data[23] ;
 wire \spi_sram_master_inst.data[24] ;
 wire \spi_sram_master_inst.data[25] ;
 wire \spi_sram_master_inst.data[26] ;
 wire \spi_sram_master_inst.data[27] ;
 wire \spi_sram_master_inst.data[28] ;
 wire \spi_sram_master_inst.data[29] ;
 wire \spi_sram_master_inst.data[30] ;
 wire \spi_sram_master_inst.data[31] ;
 wire \spi_sram_master_inst.data[32] ;
 wire \spi_sram_master_inst.data[33] ;
 wire \spi_sram_master_inst.data[34] ;
 wire \spi_sram_master_inst.data[35] ;
 wire \spi_sram_master_inst.data[36] ;
 wire \spi_sram_master_inst.data[37] ;
 wire \spi_sram_master_inst.data[38] ;
 wire \spi_sram_master_inst.data[39] ;
 wire \spi_sram_master_inst.data[8] ;
 wire \spi_sram_master_inst.data[9] ;
 wire \spi_sram_master_inst.dout ;
 wire \spi_sram_master_inst.state[0] ;
 wire \spi_sram_master_inst.state[1] ;
 wire \spi_sram_master_inst.state[2] ;
 wire \spi_sram_master_inst.state[3] ;
 wire net120;
 wire net121;
 wire net102;
 wire net122;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;

 sky130_fd_sc_hd__inv_2 _1074_ (.A(\spi_sram_master_inst.state[0] ),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(\cpu_inst.NMI_edge ),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(\cpu_inst.I ),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(net87),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _1078_ (.A(\cpu_inst.state[4] ),
    .Y(_0497_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(\cpu_inst.clc ),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(\cpu_inst.plp ),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(\cpu_inst.src_reg[1] ),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(\cpu_inst.AXYS[1][0] ),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(\cpu_inst.rotate ),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(\cpu_inst.cli ),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(\cpu_inst.cld ),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _1086_ (.A(\cpu_inst.php ),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _2148__2 (.A(clknet_4_5_0_clk),
    .Y(net123));
 sky130_fd_sc_hd__and2b_1 _1088_ (.A_N(\spi_sram_master_inst.state[3] ),
    .B(\spi_sram_master_inst.state[2] ),
    .X(_0506_));
 sky130_fd_sc_hd__nand2b_1 _1089_ (.A_N(\spi_sram_master_inst.state[3] ),
    .B(\spi_sram_master_inst.state[2] ),
    .Y(_0507_));
 sky130_fd_sc_hd__nand2_1 _1090_ (.A(\spi_sram_master_inst.state[1] ),
    .B(_0506_),
    .Y(_0508_));
 sky130_fd_sc_hd__nor3_2 _1091_ (.A(\spi_sram_master_inst.state[2] ),
    .B(\spi_sram_master_inst.state[1] ),
    .C(\spi_sram_master_inst.state[0] ),
    .Y(_0509_));
 sky130_fd_sc_hd__or3_1 _1092_ (.A(\spi_sram_master_inst.state[2] ),
    .B(\spi_sram_master_inst.state[1] ),
    .C(\spi_sram_master_inst.state[0] ),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(_0508_),
    .B(_0510_),
    .Y(\spi_sram_master_inst.cs_n_sm ));
 sky130_fd_sc_hd__or3_2 _1094_ (.A(\spi_sram_master_inst.state[1] ),
    .B(_0493_),
    .C(_0507_),
    .X(_0511_));
 sky130_fd_sc_hd__or3b_1 _1095_ (.A(\spi_sram_master_inst.state[3] ),
    .B(\spi_sram_master_inst.state[2] ),
    .C_N(\spi_sram_master_inst.state[1] ),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _1096_ (.A(_0493_),
    .B(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _1097_ (.A(_0510_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__or2_1 _1098_ (.A(\spi_sram_master_inst.counter[0] ),
    .B(\spi_sram_master_inst.counter[1] ),
    .X(_0515_));
 sky130_fd_sc_hd__xnor2_1 _1099_ (.A(\spi_sram_master_inst.counter[2] ),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__o21a_1 _1100_ (.A1(_0514_),
    .A2(_0516_),
    .B1(_0511_),
    .X(_0001_));
 sky130_fd_sc_hd__or3_1 _1101_ (.A(\spi_sram_master_inst.counter[3] ),
    .B(\spi_sram_master_inst.counter[2] ),
    .C(_0515_),
    .X(_0517_));
 sky130_fd_sc_hd__o21ai_1 _1102_ (.A1(\spi_sram_master_inst.counter[2] ),
    .A2(_0515_),
    .B1(\spi_sram_master_inst.counter[3] ),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _1103_ (.A(_0517_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_2 _1104_ (.A(_0511_),
    .B(_0513_),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _1105_ (.A(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__a31o_1 _1106_ (.A1(_0511_),
    .A2(_0513_),
    .A3(_0519_),
    .B1(_0509_),
    .X(_0002_));
 sky130_fd_sc_hd__or2_1 _1107_ (.A(_0509_),
    .B(_0520_),
    .X(_0522_));
 sky130_fd_sc_hd__nor3_1 _1108_ (.A(net128),
    .B(_0517_),
    .C(_0522_),
    .Y(_0185_));
 sky130_fd_sc_hd__a311o_1 _1109_ (.A1(net128),
    .A2(_0517_),
    .A3(_0521_),
    .B1(_0185_),
    .C1(_0509_),
    .X(_0003_));
 sky130_fd_sc_hd__o21a_1 _1110_ (.A1(\spi_sram_master_inst.state[1] ),
    .A2(_0507_),
    .B1(_0512_),
    .X(_0523_));
 sky130_fd_sc_hd__o21ai_2 _1111_ (.A1(\spi_sram_master_inst.state[1] ),
    .A2(_0507_),
    .B1(_0512_),
    .Y(_0524_));
 sky130_fd_sc_hd__mux2_1 _1112_ (.A0(_0508_),
    .A1(net70),
    .S(_0493_),
    .X(_0525_));
 sky130_fd_sc_hd__inv_2 _1113_ (.A(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__a211oi_1 _1114_ (.A1(\spi_sram_master_inst.state[3] ),
    .A2(_0509_),
    .B1(_0520_),
    .C1(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__a211o_2 _1115_ (.A1(\spi_sram_master_inst.state[3] ),
    .A2(_0509_),
    .B1(_0520_),
    .C1(_0526_),
    .X(_0528_));
 sky130_fd_sc_hd__and2b_1 _1116_ (.A_N(\cpu_inst.state[5] ),
    .B(\cpu_inst.state[4] ),
    .X(_0529_));
 sky130_fd_sc_hd__nand2b_1 _1117_ (.A_N(\cpu_inst.state[5] ),
    .B(\cpu_inst.state[4] ),
    .Y(_0530_));
 sky130_fd_sc_hd__and4b_1 _1118_ (.A_N(net90),
    .B(net92),
    .C(net86),
    .D(net88),
    .X(_0531_));
 sky130_fd_sc_hd__or4bb_1 _1119_ (.A(_0496_),
    .B(net91),
    .C_N(net93),
    .D_N(net89),
    .X(_0532_));
 sky130_fd_sc_hd__and2b_1 _1120_ (.A_N(\cpu_inst.state[4] ),
    .B(\cpu_inst.state[5] ),
    .X(_0533_));
 sky130_fd_sc_hd__nand2b_2 _1121_ (.A_N(\cpu_inst.state[4] ),
    .B(\cpu_inst.state[5] ),
    .Y(_0534_));
 sky130_fd_sc_hd__o21a_1 _1122_ (.A1(_0529_),
    .A2(_0533_),
    .B1(_0531_),
    .X(_0535_));
 sky130_fd_sc_hd__and4b_1 _1123_ (.A_N(net92),
    .B(net86),
    .C(net88),
    .D(net90),
    .X(_0536_));
 sky130_fd_sc_hd__and2_1 _1124_ (.A(_0533_),
    .B(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__or4b_4 _1125_ (.A(net91),
    .B(net87),
    .C(net89),
    .D_N(net92),
    .X(_0538_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__nor2_1 _1127_ (.A(net76),
    .B(_0538_),
    .Y(_0540_));
 sky130_fd_sc_hd__and2b_1 _1128_ (.A_N(net87),
    .B(net88),
    .X(_0541_));
 sky130_fd_sc_hd__or4bb_2 _1129_ (.A(net91),
    .B(net86),
    .C_N(net89),
    .D_N(net92),
    .X(_0542_));
 sky130_fd_sc_hd__nor2_1 _1130_ (.A(net75),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__or4_1 _1131_ (.A(_0535_),
    .B(net66),
    .C(_0540_),
    .D(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__or3b_4 _1132_ (.A(net91),
    .B(net93),
    .C_N(_0541_),
    .X(_0545_));
 sky130_fd_sc_hd__nor2_1 _1133_ (.A(net75),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__or2_1 _1134_ (.A(\cpu_inst.ALU.CO ),
    .B(\cpu_inst.store ),
    .X(_0547_));
 sky130_fd_sc_hd__or3_1 _1135_ (.A(net76),
    .B(_0545_),
    .C(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__and2_1 _1136_ (.A(net91),
    .B(net93),
    .X(_0549_));
 sky130_fd_sc_hd__nand4_2 _1137_ (.A(net90),
    .B(net92),
    .C(net86),
    .D(net88),
    .Y(_0550_));
 sky130_fd_sc_hd__nor2_1 _1138_ (.A(net74),
    .B(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__nor2_1 _1139_ (.A(\cpu_inst.state[5] ),
    .B(\cpu_inst.state[4] ),
    .Y(_0552_));
 sky130_fd_sc_hd__or2_1 _1140_ (.A(\cpu_inst.state[5] ),
    .B(\cpu_inst.state[4] ),
    .X(_0553_));
 sky130_fd_sc_hd__nor2_1 _1141_ (.A(_0545_),
    .B(net73),
    .Y(_0554_));
 sky130_fd_sc_hd__or2_1 _1142_ (.A(_0551_),
    .B(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _1143_ (.A(_0538_),
    .B(net73),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _1144_ (.A(\cpu_inst.state[5] ),
    .B(\cpu_inst.state[4] ),
    .Y(_0557_));
 sky130_fd_sc_hd__nor2_1 _1145_ (.A(_0538_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__or3_1 _1146_ (.A(_0555_),
    .B(_0556_),
    .C(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__or4bb_2 _1147_ (.A(net86),
    .B(net88),
    .C_N(net90),
    .D_N(net92),
    .X(_0560_));
 sky130_fd_sc_hd__nor2_2 _1148_ (.A(net72),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__o21ba_1 _1149_ (.A1(_0546_),
    .A2(_0561_),
    .B1_N(_0547_),
    .X(_0562_));
 sky130_fd_sc_hd__o2bb2a_1 _1150_ (.A1_N(\cpu_inst.write_back ),
    .A2_N(_0548_),
    .B1(_0559_),
    .B2(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__or4bb_2 _1151_ (.A(net90),
    .B(net92),
    .C_N(net86),
    .D_N(net88),
    .X(_0564_));
 sky130_fd_sc_hd__nor2_2 _1152_ (.A(net75),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__and3_1 _1153_ (.A(net31),
    .B(_0529_),
    .C(_0531_),
    .X(_0566_));
 sky130_fd_sc_hd__a21o_1 _1154_ (.A1(net38),
    .A2(_0565_),
    .B1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_4 _1155_ (.A(_0532_),
    .B(net73),
    .Y(_0568_));
 sky130_fd_sc_hd__nor2_1 _1156_ (.A(net74),
    .B(_0564_),
    .Y(_0569_));
 sky130_fd_sc_hd__and3_1 _1157_ (.A(net31),
    .B(_0531_),
    .C(_0533_),
    .X(_0570_));
 sky130_fd_sc_hd__a21o_1 _1158_ (.A1(net38),
    .A2(_0569_),
    .B1(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__nor2_1 _1159_ (.A(net72),
    .B(_0564_),
    .Y(_0572_));
 sky130_fd_sc_hd__or2_4 _1160_ (.A(net72),
    .B(_0564_),
    .X(_0573_));
 sky130_fd_sc_hd__nor2_1 _1161_ (.A(net29),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_1 _1162_ (.A(net36),
    .B(net65),
    .Y(_0575_));
 sky130_fd_sc_hd__and2b_1 _1163_ (.A_N(net77),
    .B(\cpu_inst.DI[4] ),
    .X(_0576_));
 sky130_fd_sc_hd__a21oi_2 _1164_ (.A1(net77),
    .A2(\cpu_inst.IRHOLD[4] ),
    .B1(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__a21o_2 _1165_ (.A1(net77),
    .A2(\cpu_inst.IRHOLD[4] ),
    .B1(_0576_),
    .X(_0578_));
 sky130_fd_sc_hd__a21oi_1 _1166_ (.A1(_0495_),
    .A2(net2),
    .B1(\cpu_inst.NMI_edge ),
    .Y(_0579_));
 sky130_fd_sc_hd__and2_1 _1167_ (.A(_0578_),
    .B(net62),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_1 _1168_ (.A(_0578_),
    .B(net62),
    .Y(_0581_));
 sky130_fd_sc_hd__mux2_2 _1169_ (.A0(net97),
    .A1(\cpu_inst.IRHOLD[2] ),
    .S(net77),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _1170_ (.A0(net96),
    .A1(\cpu_inst.IRHOLD[3] ),
    .S(net77),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _1171_ (.A(net62),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__or2_2 _1172_ (.A(_0582_),
    .B(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_2 _1173_ (.A0(net99),
    .A1(\cpu_inst.IRHOLD[0] ),
    .S(net77),
    .X(_0586_));
 sky130_fd_sc_hd__nand2_1 _1174_ (.A(net62),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(net98),
    .A1(\cpu_inst.IRHOLD[1] ),
    .S(net77),
    .X(_0588_));
 sky130_fd_sc_hd__or2_4 _1176_ (.A(_0587_),
    .B(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__inv_2 _1177_ (.A(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nor2_1 _1178_ (.A(_0585_),
    .B(_0589_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _1179_ (.A(net62),
    .B(_0582_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(_0584_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__mux2_4 _1181_ (.A0(net94),
    .A1(\cpu_inst.IRHOLD[7] ),
    .S(net77),
    .X(_0594_));
 sky130_fd_sc_hd__and2_2 _1182_ (.A(net63),
    .B(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_4 _1183_ (.A(net63),
    .B(_0594_),
    .Y(_0596_));
 sky130_fd_sc_hd__o32a_1 _1184_ (.A1(_0586_),
    .A2(_0593_),
    .A3(_0596_),
    .B1(_0589_),
    .B2(_0585_),
    .X(_0597_));
 sky130_fd_sc_hd__nor2_1 _1185_ (.A(net50),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__a211o_1 _1186_ (.A1(net65),
    .A2(_0598_),
    .B1(_0544_),
    .C1(_0563_),
    .X(_0599_));
 sky130_fd_sc_hd__a211o_1 _1187_ (.A1(net37),
    .A2(_0599_),
    .B1(_0571_),
    .C1(_0567_),
    .X(_0600_));
 sky130_fd_sc_hd__a21o_1 _1188_ (.A1(net29),
    .A2(_0568_),
    .B1(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__nand2_2 _1189_ (.A(net62),
    .B(_0588_),
    .Y(_0602_));
 sky130_fd_sc_hd__inv_2 _1190_ (.A(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__and2_1 _1191_ (.A(_0587_),
    .B(_0602_),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_1 _1192_ (.A(_0587_),
    .B(_0602_),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _1193_ (.A(_0593_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__mux2_2 _1194_ (.A0(\cpu_inst.DI[5] ),
    .A1(\cpu_inst.IRHOLD[5] ),
    .S(net77),
    .X(_0607_));
 sky130_fd_sc_hd__inv_2 _1195_ (.A(net71),
    .Y(_0608_));
 sky130_fd_sc_hd__nor2_1 _1196_ (.A(_0578_),
    .B(net71),
    .Y(_0609_));
 sky130_fd_sc_hd__and2_2 _1197_ (.A(net63),
    .B(_0607_),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_1 _1198_ (.A(net62),
    .B(net71),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _1199_ (.A(net50),
    .B(_0610_),
    .Y(_0612_));
 sky130_fd_sc_hd__mux2_2 _1200_ (.A0(net95),
    .A1(\cpu_inst.IRHOLD[6] ),
    .S(\cpu_inst.IRHOLD_valid ),
    .X(_0613_));
 sky130_fd_sc_hd__and2_1 _1201_ (.A(net63),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__nand2_2 _1202_ (.A(net63),
    .B(_0613_),
    .Y(_0615_));
 sky130_fd_sc_hd__or2_1 _1203_ (.A(_0594_),
    .B(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__inv_2 _1204_ (.A(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _1205_ (.A(net19),
    .B(_0616_),
    .Y(_0618_));
 sky130_fd_sc_hd__nor2_2 _1206_ (.A(net74),
    .B(_0542_),
    .Y(_0619_));
 sky130_fd_sc_hd__a32o_1 _1207_ (.A1(_0606_),
    .A2(_0612_),
    .A3(_0618_),
    .B1(_0619_),
    .B2(net29),
    .X(_0620_));
 sky130_fd_sc_hd__nor2_2 _1208_ (.A(_0542_),
    .B(net72),
    .Y(_0621_));
 sky130_fd_sc_hd__a32o_1 _1209_ (.A1(net21),
    .A2(net50),
    .A3(_0606_),
    .B1(net61),
    .B2(net29),
    .X(_0622_));
 sky130_fd_sc_hd__and3_1 _1210_ (.A(net39),
    .B(_0546_),
    .C(_0547_),
    .X(_0623_));
 sky130_fd_sc_hd__a21o_1 _1211_ (.A1(net31),
    .A2(_0543_),
    .B1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or4_1 _1212_ (.A(_0601_),
    .B(_0620_),
    .C(_0622_),
    .D(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__and2_1 _1213_ (.A(net31),
    .B(_0551_),
    .X(_0626_));
 sky130_fd_sc_hd__nor2_1 _1214_ (.A(_0583_),
    .B(_0592_),
    .Y(_0627_));
 sky130_fd_sc_hd__or3b_1 _1215_ (.A(net19),
    .B(_0578_),
    .C_N(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__nor2_1 _1216_ (.A(_0550_),
    .B(net72),
    .Y(_0629_));
 sky130_fd_sc_hd__and2_1 _1217_ (.A(_0536_),
    .B(_0552_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _1218_ (.A0(_0629_),
    .A1(_0630_),
    .S(net36),
    .X(_0631_));
 sky130_fd_sc_hd__or3b_1 _1219_ (.A(_0626_),
    .B(_0631_),
    .C_N(_0628_),
    .X(_0632_));
 sky130_fd_sc_hd__or4bb_2 _1220_ (.A(net92),
    .B(net86),
    .C_N(net88),
    .D_N(net90),
    .X(_0633_));
 sky130_fd_sc_hd__nor2_1 _1221_ (.A(net75),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__and3_2 _1222_ (.A(_0529_),
    .B(_0541_),
    .C(_0549_),
    .X(_0635_));
 sky130_fd_sc_hd__nor2_1 _1223_ (.A(net75),
    .B(_0550_),
    .Y(_0636_));
 sky130_fd_sc_hd__or2_1 _1224_ (.A(net38),
    .B(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__and2_2 _1225_ (.A(_0529_),
    .B(_0536_),
    .X(_0638_));
 sky130_fd_sc_hd__o21ai_1 _1226_ (.A1(net28),
    .A2(_0638_),
    .B1(_0637_),
    .Y(_0639_));
 sky130_fd_sc_hd__a21bo_1 _1227_ (.A1(net30),
    .A2(_0635_),
    .B1_N(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__a21o_1 _1228_ (.A1(net36),
    .A2(_0634_),
    .B1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__and3_2 _1229_ (.A(_0541_),
    .B(_0549_),
    .C(_0552_),
    .X(_0642_));
 sky130_fd_sc_hd__nor2_1 _1230_ (.A(net73),
    .B(_0633_),
    .Y(_0643_));
 sky130_fd_sc_hd__xnor2_2 _1231_ (.A(\cpu_inst.backwards ),
    .B(\cpu_inst.ALU.CO ),
    .Y(_0644_));
 sky130_fd_sc_hd__inv_2 _1232_ (.A(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__and3_1 _1233_ (.A(net37),
    .B(net55),
    .C(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__and3_1 _1234_ (.A(_0533_),
    .B(_0541_),
    .C(_0549_),
    .X(_0647_));
 sky130_fd_sc_hd__nor2_1 _1235_ (.A(net74),
    .B(_0633_),
    .Y(_0648_));
 sky130_fd_sc_hd__mux2_1 _1236_ (.A0(net54),
    .A1(_0648_),
    .S(net37),
    .X(_0649_));
 sky130_fd_sc_hd__a211o_1 _1237_ (.A1(_0528_),
    .A2(net60),
    .B1(_0646_),
    .C1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__or3_1 _1238_ (.A(_0632_),
    .B(_0641_),
    .C(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__and2b_1 _1239_ (.A_N(net89),
    .B(net87),
    .X(_0652_));
 sky130_fd_sc_hd__or4b_2 _1240_ (.A(net91),
    .B(net89),
    .C(_0496_),
    .D_N(net93),
    .X(_0653_));
 sky130_fd_sc_hd__nor2_1 _1241_ (.A(_0534_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__or4b_4 _1242_ (.A(net90),
    .B(net93),
    .C(net89),
    .D_N(net87),
    .X(_0655_));
 sky130_fd_sc_hd__nor2_1 _1243_ (.A(\cpu_inst.state[4] ),
    .B(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__nor2_1 _1244_ (.A(net74),
    .B(_0655_),
    .Y(_0657_));
 sky130_fd_sc_hd__mux2_1 _1245_ (.A0(_0654_),
    .A1(_0657_),
    .S(net38),
    .X(_0658_));
 sky130_fd_sc_hd__nor2_1 _1246_ (.A(net75),
    .B(_0653_),
    .Y(_0659_));
 sky130_fd_sc_hd__nor2_1 _1247_ (.A(net75),
    .B(_0655_),
    .Y(_0660_));
 sky130_fd_sc_hd__mux2_1 _1248_ (.A0(_0659_),
    .A1(_0660_),
    .S(net36),
    .X(_0661_));
 sky130_fd_sc_hd__nor2_1 _1249_ (.A(net73),
    .B(_0655_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand2_1 _1250_ (.A(net39),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__inv_2 _1251_ (.A(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__nor2_2 _1252_ (.A(net72),
    .B(_0653_),
    .Y(_0665_));
 sky130_fd_sc_hd__a2111o_1 _1253_ (.A1(net28),
    .A2(_0665_),
    .B1(_0664_),
    .C1(_0661_),
    .D1(_0658_),
    .X(_0666_));
 sky130_fd_sc_hd__or4_4 _1254_ (.A(net90),
    .B(net92),
    .C(net86),
    .D(net88),
    .X(_0667_));
 sky130_fd_sc_hd__nor2_1 _1255_ (.A(_0557_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__mux2_1 _1256_ (.A0(_0558_),
    .A1(_0668_),
    .S(net38),
    .X(_0669_));
 sky130_fd_sc_hd__nor2_1 _1257_ (.A(\cpu_inst.state[5] ),
    .B(_0667_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _1258_ (.A(net75),
    .B(_0667_),
    .Y(_0671_));
 sky130_fd_sc_hd__mux2_1 _1259_ (.A0(_0540_),
    .A1(_0671_),
    .S(net40),
    .X(_0672_));
 sky130_fd_sc_hd__or2_1 _1260_ (.A(_0669_),
    .B(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_1 _1261_ (.A(net72),
    .B(_0667_),
    .Y(_0674_));
 sky130_fd_sc_hd__mux2_1 _1262_ (.A0(_0556_),
    .A1(_0674_),
    .S(net37),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_2 _1263_ (.A(_0585_),
    .B(_0605_),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_1 _1264_ (.A(_0612_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nor2_1 _1265_ (.A(_0595_),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__and2_1 _1266_ (.A(net20),
    .B(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__nor2_1 _1267_ (.A(net74),
    .B(_0538_),
    .Y(_0680_));
 sky130_fd_sc_hd__a2111o_1 _1268_ (.A1(net29),
    .A2(_0680_),
    .B1(_0679_),
    .C1(_0675_),
    .D1(_0673_),
    .X(_0681_));
 sky130_fd_sc_hd__and3_2 _1269_ (.A(_0549_),
    .B(_0552_),
    .C(_0652_),
    .X(_0682_));
 sky130_fd_sc_hd__or4bb_4 _1270_ (.A(net93),
    .B(net89),
    .C_N(net87),
    .D_N(net91),
    .X(_0683_));
 sky130_fd_sc_hd__nor2_1 _1271_ (.A(\cpu_inst.state[5] ),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__nor2_2 _1272_ (.A(net73),
    .B(_0683_),
    .Y(_0685_));
 sky130_fd_sc_hd__or2_1 _1273_ (.A(net73),
    .B(_0683_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(_0682_),
    .A1(net52),
    .S(net37),
    .X(_0687_));
 sky130_fd_sc_hd__and3_1 _1275_ (.A(_0533_),
    .B(_0549_),
    .C(_0652_),
    .X(_0688_));
 sky130_fd_sc_hd__or2_1 _1276_ (.A(net38),
    .B(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__nor2_1 _1277_ (.A(net74),
    .B(_0683_),
    .Y(_0690_));
 sky130_fd_sc_hd__o21ai_1 _1278_ (.A1(net29),
    .A2(_0690_),
    .B1(_0689_),
    .Y(_0691_));
 sky130_fd_sc_hd__inv_2 _1279_ (.A(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2_4 _1280_ (.A(net76),
    .B(_0683_),
    .Y(_0693_));
 sky130_fd_sc_hd__or2_4 _1281_ (.A(net76),
    .B(_0683_),
    .X(_0694_));
 sky130_fd_sc_hd__and3_2 _1282_ (.A(_0529_),
    .B(_0549_),
    .C(_0652_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _1283_ (.A0(_0693_),
    .A1(_0695_),
    .S(net28),
    .X(_0696_));
 sky130_fd_sc_hd__or3_1 _1284_ (.A(_0687_),
    .B(_0692_),
    .C(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__nor2_2 _1285_ (.A(net75),
    .B(_0560_),
    .Y(_0698_));
 sky130_fd_sc_hd__or4b_4 _1286_ (.A(net92),
    .B(net86),
    .C(net88),
    .D_N(net90),
    .X(_0699_));
 sky130_fd_sc_hd__nor2_2 _1287_ (.A(net75),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__mux2_1 _1288_ (.A0(_0698_),
    .A1(_0700_),
    .S(net36),
    .X(_0701_));
 sky130_fd_sc_hd__and3_1 _1289_ (.A(\cpu_inst.write_back ),
    .B(net39),
    .C(_0559_),
    .X(_0702_));
 sky130_fd_sc_hd__nor2_2 _1290_ (.A(net74),
    .B(_0560_),
    .Y(_0703_));
 sky130_fd_sc_hd__a21o_1 _1291_ (.A1(net31),
    .A2(_0703_),
    .B1(_0702_),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_2 _1292_ (.A(net72),
    .B(_0699_),
    .Y(_0705_));
 sky130_fd_sc_hd__mux2_1 _1293_ (.A0(_0561_),
    .A1(_0705_),
    .S(net36),
    .X(_0706_));
 sky130_fd_sc_hd__or3_1 _1294_ (.A(_0701_),
    .B(_0704_),
    .C(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__or3_1 _1295_ (.A(_0651_),
    .B(_0697_),
    .C(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__or4_1 _1296_ (.A(_0625_),
    .B(_0666_),
    .C(_0681_),
    .D(_0708_),
    .X(_0004_));
 sky130_fd_sc_hd__nor2_1 _1297_ (.A(_0589_),
    .B(_0593_),
    .Y(_0709_));
 sky130_fd_sc_hd__a32o_1 _1298_ (.A1(net20),
    .A2(net50),
    .A3(_0709_),
    .B1(_0700_),
    .B2(net28),
    .X(_0710_));
 sky130_fd_sc_hd__and3_1 _1299_ (.A(net62),
    .B(_0582_),
    .C(_0583_),
    .X(_0711_));
 sky130_fd_sc_hd__o21a_1 _1300_ (.A1(_0591_),
    .A2(_0711_),
    .B1(net50),
    .X(_0712_));
 sky130_fd_sc_hd__or2_1 _1301_ (.A(net30),
    .B(_0665_),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _1302_ (.A1(net20),
    .A2(_0712_),
    .B1(_0713_),
    .B2(_0705_),
    .X(_0714_));
 sky130_fd_sc_hd__o21a_1 _1303_ (.A1(net36),
    .A2(net52),
    .B1(_0713_),
    .X(_0715_));
 sky130_fd_sc_hd__nor2_4 _1304_ (.A(net74),
    .B(_0699_),
    .Y(_0716_));
 sky130_fd_sc_hd__mux2_1 _1305_ (.A0(_0680_),
    .A1(_0716_),
    .S(net30),
    .X(_0717_));
 sky130_fd_sc_hd__or4_1 _1306_ (.A(_0710_),
    .B(_0714_),
    .C(_0715_),
    .D(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__nor2_1 _1307_ (.A(_0578_),
    .B(_0611_),
    .Y(_0719_));
 sky130_fd_sc_hd__and3_1 _1308_ (.A(_0606_),
    .B(_0617_),
    .C(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__a22o_1 _1309_ (.A1(net29),
    .A2(_0690_),
    .B1(_0720_),
    .B2(net21),
    .X(_0721_));
 sky130_fd_sc_hd__and3_1 _1310_ (.A(_0596_),
    .B(_0615_),
    .C(_0719_),
    .X(_0722_));
 sky130_fd_sc_hd__and2_1 _1311_ (.A(_0606_),
    .B(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__a22o_1 _1312_ (.A1(net28),
    .A2(_0693_),
    .B1(_0723_),
    .B2(net20),
    .X(_0724_));
 sky130_fd_sc_hd__or2_1 _1313_ (.A(_0721_),
    .B(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__and3_1 _1314_ (.A(_0596_),
    .B(_0676_),
    .C(_0719_),
    .X(_0726_));
 sky130_fd_sc_hd__and2_1 _1315_ (.A(net21),
    .B(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__a21o_1 _1316_ (.A1(net28),
    .A2(_0638_),
    .B1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _1317_ (.A0(net66),
    .A1(_0703_),
    .S(net36),
    .X(_0729_));
 sky130_fd_sc_hd__a32o_1 _1318_ (.A1(net20),
    .A2(_0581_),
    .A3(_0709_),
    .B1(_0630_),
    .B2(net28),
    .X(_0730_));
 sky130_fd_sc_hd__or3_1 _1319_ (.A(_0728_),
    .B(_0729_),
    .C(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__and3_1 _1320_ (.A(_0587_),
    .B(_0602_),
    .C(_0711_),
    .X(_0732_));
 sky130_fd_sc_hd__and3_1 _1321_ (.A(_0609_),
    .B(_0617_),
    .C(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__o21a_1 _1322_ (.A1(_0659_),
    .A2(_0682_),
    .B1(net36),
    .X(_0734_));
 sky130_fd_sc_hd__a221o_1 _1323_ (.A1(net28),
    .A2(_0634_),
    .B1(_0733_),
    .B2(net21),
    .C1(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(_0619_),
    .A1(_0648_),
    .S(net31),
    .X(_0736_));
 sky130_fd_sc_hd__mux4_2 _1325_ (.A0(\cpu_inst.N ),
    .A1(\cpu_inst.V ),
    .A2(\cpu_inst.C ),
    .A3(\cpu_inst.Z ),
    .S0(\cpu_inst.cond_code[1] ),
    .S1(\cpu_inst.cond_code[2] ),
    .X(_0737_));
 sky130_fd_sc_hd__xnor2_1 _1326_ (.A(\cpu_inst.cond_code[0] ),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__and3_1 _1327_ (.A(net37),
    .B(net61),
    .C(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__a211o_1 _1328_ (.A1(_0528_),
    .A2(net55),
    .B1(_0736_),
    .C1(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__or3_1 _1329_ (.A(_0731_),
    .B(_0735_),
    .C(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__or4_1 _1330_ (.A(_0708_),
    .B(_0718_),
    .C(_0725_),
    .D(_0741_),
    .X(_0005_));
 sky130_fd_sc_hd__and3_1 _1331_ (.A(_0596_),
    .B(_0606_),
    .C(_0612_),
    .X(_0742_));
 sky130_fd_sc_hd__a21o_1 _1332_ (.A1(_0577_),
    .A2(_0595_),
    .B1(_0722_),
    .X(_0743_));
 sky130_fd_sc_hd__nor2_1 _1333_ (.A(_0586_),
    .B(_0602_),
    .Y(_0744_));
 sky130_fd_sc_hd__or2_2 _1334_ (.A(_0586_),
    .B(_0602_),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_1 _1335_ (.A(_0589_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__a32o_1 _1336_ (.A1(_0577_),
    .A2(_0711_),
    .A3(_0746_),
    .B1(_0743_),
    .B2(_0732_),
    .X(_0747_));
 sky130_fd_sc_hd__a211o_1 _1337_ (.A1(net50),
    .A2(_0606_),
    .B1(_0627_),
    .C1(_0709_),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_1 _1338_ (.A(_0585_),
    .B(_0586_),
    .Y(_0749_));
 sky130_fd_sc_hd__o31a_1 _1339_ (.A1(_0578_),
    .A2(_0595_),
    .A3(_0603_),
    .B1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__and3_1 _1340_ (.A(_0617_),
    .B(_0719_),
    .C(_0732_),
    .X(_0751_));
 sky130_fd_sc_hd__or4_1 _1341_ (.A(_0678_),
    .B(_0720_),
    .C(_0723_),
    .D(_0748_),
    .X(_0752_));
 sky130_fd_sc_hd__or4_1 _1342_ (.A(_0598_),
    .B(_0726_),
    .C(_0742_),
    .D(_0750_),
    .X(_0753_));
 sky130_fd_sc_hd__or4_1 _1343_ (.A(_0712_),
    .B(_0733_),
    .C(_0751_),
    .D(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__o31a_1 _1344_ (.A1(_0747_),
    .A2(_0752_),
    .A3(_0754_),
    .B1(net37),
    .X(_0755_));
 sky130_fd_sc_hd__nor2_1 _1345_ (.A(_0573_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__a2111o_1 _1346_ (.A1(net55),
    .A2(_0644_),
    .B1(_0568_),
    .C1(_0635_),
    .D1(net60),
    .X(_0757_));
 sky130_fd_sc_hd__nor2_1 _1347_ (.A(net74),
    .B(_0667_),
    .Y(_0758_));
 sky130_fd_sc_hd__nor2_4 _1348_ (.A(_0534_),
    .B(_0545_),
    .Y(_0759_));
 sky130_fd_sc_hd__or4_1 _1349_ (.A(_0654_),
    .B(_0716_),
    .C(_0758_),
    .D(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__nor2_1 _1350_ (.A(_0757_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__o31ai_1 _1351_ (.A1(_0542_),
    .A2(net72),
    .A3(_0738_),
    .B1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__mux2_1 _1352_ (.A0(_0565_),
    .A1(_0695_),
    .S(net36),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _1353_ (.A0(_0569_),
    .A1(_0688_),
    .S(net38),
    .X(_0764_));
 sky130_fd_sc_hd__a2111o_1 _1354_ (.A1(net37),
    .A2(_0762_),
    .B1(_0763_),
    .C1(_0764_),
    .D1(_0756_),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _1355_ (.A1(net21),
    .A2(_0750_),
    .B1(_0759_),
    .B2(net29),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(_0546_),
    .A1(_0698_),
    .S(net39),
    .X(_0767_));
 sky130_fd_sc_hd__o211a_1 _1357_ (.A1(\cpu_inst.write_back ),
    .A2(_0547_),
    .B1(_0561_),
    .C1(net39),
    .X(_0768_));
 sky130_fd_sc_hd__a211o_1 _1358_ (.A1(net31),
    .A2(_0554_),
    .B1(_0767_),
    .C1(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__or4_1 _1359_ (.A(_0741_),
    .B(_0765_),
    .C(_0766_),
    .D(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__or3_1 _1360_ (.A(_0625_),
    .B(_0651_),
    .C(_0770_),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _1361_ (.A1(net28),
    .A2(_0660_),
    .B1(_0751_),
    .B2(net21),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(net54),
    .A1(_0657_),
    .S(net29),
    .X(_0772_));
 sky130_fd_sc_hd__or3_1 _1363_ (.A(_0725_),
    .B(_0771_),
    .C(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__a32o_1 _1364_ (.A1(net21),
    .A2(_0578_),
    .A3(_0627_),
    .B1(_0668_),
    .B2(net28),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _1365_ (.A0(_0629_),
    .A1(_0671_),
    .S(net30),
    .X(_0775_));
 sky130_fd_sc_hd__or2_1 _1366_ (.A(_0774_),
    .B(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__or2_2 _1367_ (.A(net30),
    .B(_0636_),
    .X(_0777_));
 sky130_fd_sc_hd__o21a_1 _1368_ (.A1(net37),
    .A2(_0758_),
    .B1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__a221o_1 _1369_ (.A1(net20),
    .A2(_0747_),
    .B1(_0777_),
    .B2(_0674_),
    .C1(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__or4_1 _1370_ (.A(_0718_),
    .B(_0773_),
    .C(_0776_),
    .D(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__or3_1 _1371_ (.A(_0004_),
    .B(_0770_),
    .C(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__or4b_1 _1372_ (.A(_0632_),
    .B(_0731_),
    .C(_0715_),
    .D_N(_0639_),
    .X(_0782_));
 sky130_fd_sc_hd__or4_1 _1373_ (.A(_0666_),
    .B(_0697_),
    .C(_0773_),
    .D(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__or4b_1 _1374_ (.A(_0601_),
    .B(_0765_),
    .C(_0783_),
    .D_N(_0781_),
    .X(_0007_));
 sky130_fd_sc_hd__or3_1 _1375_ (.A(_0724_),
    .B(_0728_),
    .C(_0771_),
    .X(_0784_));
 sky130_fd_sc_hd__or4_1 _1376_ (.A(_0661_),
    .B(_0710_),
    .C(_0763_),
    .D(_0767_),
    .X(_0785_));
 sky130_fd_sc_hd__or4_1 _1377_ (.A(_0567_),
    .B(_0624_),
    .C(_0673_),
    .D(_0696_),
    .X(_0786_));
 sky130_fd_sc_hd__or4_1 _1378_ (.A(_0641_),
    .B(_0701_),
    .C(_0785_),
    .D(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__or4_1 _1379_ (.A(_0735_),
    .B(_0776_),
    .C(_0784_),
    .D(_0787_),
    .X(_0008_));
 sky130_fd_sc_hd__or4_1 _1380_ (.A(_0736_),
    .B(_0764_),
    .C(_0772_),
    .D(_0778_),
    .X(_0788_));
 sky130_fd_sc_hd__or3b_1 _1381_ (.A(_0626_),
    .B(_0774_),
    .C_N(_0628_),
    .X(_0789_));
 sky130_fd_sc_hd__a211o_1 _1382_ (.A1(net29),
    .A2(_0680_),
    .B1(_0721_),
    .C1(_0679_),
    .X(_0790_));
 sky130_fd_sc_hd__or4_1 _1383_ (.A(_0658_),
    .B(_0669_),
    .C(_0717_),
    .D(_0729_),
    .X(_0791_));
 sky130_fd_sc_hd__or4_1 _1384_ (.A(_0571_),
    .B(_0649_),
    .C(_0692_),
    .D(_0704_),
    .X(_0792_));
 sky130_fd_sc_hd__or4_1 _1385_ (.A(_0766_),
    .B(_0790_),
    .C(_0791_),
    .D(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__or4_1 _1386_ (.A(_0620_),
    .B(_0788_),
    .C(_0789_),
    .D(_0793_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _1387_ (.A(net254),
    .B(\cpu_inst.adc_sbc ),
    .X(_0000_));
 sky130_fd_sc_hd__or3b_1 _1388_ (.A(_0509_),
    .B(_0520_),
    .C_N(net234),
    .X(_0012_));
 sky130_fd_sc_hd__nand2_1 _1389_ (.A(\spi_sram_master_inst.counter[0] ),
    .B(net196),
    .Y(_0794_));
 sky130_fd_sc_hd__a21oi_1 _1390_ (.A1(_0515_),
    .A2(net197),
    .B1(_0522_),
    .Y(_0013_));
 sky130_fd_sc_hd__and2_1 _1391_ (.A(\spi_sram_master_inst.cs_n_sm ),
    .B(net31),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_1 _1392_ (.A(\spi_sram_master_inst.cs_n_sm ),
    .B(net31),
    .Y(_0796_));
 sky130_fd_sc_hd__a21oi_2 _1393_ (.A1(net76),
    .A2(_0534_),
    .B1(_0683_),
    .Y(_0797_));
 sky130_fd_sc_hd__or4_1 _1394_ (.A(_0565_),
    .B(_0569_),
    .C(_0656_),
    .D(_0716_),
    .X(_0798_));
 sky130_fd_sc_hd__and4_1 _1395_ (.A(net90),
    .B(net86),
    .C(net88),
    .D(_0529_),
    .X(_0799_));
 sky130_fd_sc_hd__or4_1 _1396_ (.A(_0619_),
    .B(_0682_),
    .C(_0797_),
    .D(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__o22a_1 _1397_ (.A1(_0557_),
    .A2(_0667_),
    .B1(_0699_),
    .B2(net72),
    .X(_0801_));
 sky130_fd_sc_hd__or3b_2 _1398_ (.A(_0630_),
    .B(_0698_),
    .C_N(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__nor4b_1 _1399_ (.A(net65),
    .B(_0630_),
    .C(_0698_),
    .D_N(_0801_),
    .Y(_0803_));
 sky130_fd_sc_hd__or4b_2 _1400_ (.A(\cpu_inst.src_reg[0] ),
    .B(_0798_),
    .C(_0800_),
    .D_N(net48),
    .X(_0804_));
 sky130_fd_sc_hd__and2_1 _1401_ (.A(\cpu_inst.dst_reg[0] ),
    .B(net65),
    .X(_0805_));
 sky130_fd_sc_hd__a211o_1 _1402_ (.A1(\cpu_inst.index_y ),
    .A2(_0802_),
    .B1(net49),
    .C1(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(_0804_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__nor4b_1 _1404_ (.A(_0500_),
    .B(_0798_),
    .C(_0800_),
    .D_N(net48),
    .Y(_0808_));
 sky130_fd_sc_hd__a21o_1 _1405_ (.A1(\cpu_inst.dst_reg[1] ),
    .A2(net64),
    .B1(_0802_),
    .X(_0809_));
 sky130_fd_sc_hd__nor2_4 _1406_ (.A(net45),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__or2_4 _1407_ (.A(net45),
    .B(_0809_),
    .X(_0811_));
 sky130_fd_sc_hd__a21o_1 _1408_ (.A1(_0804_),
    .A2(_0806_),
    .B1(\cpu_inst.AXYS[2][0] ),
    .X(_0812_));
 sky130_fd_sc_hd__o211ai_1 _1409_ (.A1(\cpu_inst.AXYS[3][0] ),
    .A2(net26),
    .B1(_0811_),
    .C1(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand2_2 _1410_ (.A(net27),
    .B(_0810_),
    .Y(_0814_));
 sky130_fd_sc_hd__nand3_1 _1411_ (.A(\cpu_inst.AXYS[0][0] ),
    .B(net26),
    .C(_0810_),
    .Y(_0815_));
 sky130_fd_sc_hd__nor2_2 _1412_ (.A(net27),
    .B(_0811_),
    .Y(_0816_));
 sky130_fd_sc_hd__or2_2 _1413_ (.A(net26),
    .B(_0811_),
    .X(_0817_));
 sky130_fd_sc_hd__or3_1 _1414_ (.A(_0501_),
    .B(net26),
    .C(_0811_),
    .X(_0818_));
 sky130_fd_sc_hd__and3_1 _1415_ (.A(_0813_),
    .B(_0815_),
    .C(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__or2_4 _1416_ (.A(_0665_),
    .B(_0695_),
    .X(_0820_));
 sky130_fd_sc_hd__or2_2 _1417_ (.A(_0662_),
    .B(_0716_),
    .X(_0821_));
 sky130_fd_sc_hd__or3_1 _1418_ (.A(_0684_),
    .B(_0820_),
    .C(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__nor2_1 _1419_ (.A(net66),
    .B(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__nand2_4 _1420_ (.A(net40),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__nor2_1 _1421_ (.A(_0819_),
    .B(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__nor2_1 _1422_ (.A(net32),
    .B(_0823_),
    .Y(_0826_));
 sky130_fd_sc_hd__a21o_2 _1423_ (.A1(\cpu_inst.php ),
    .A2(_0716_),
    .B1(net51),
    .X(_0827_));
 sky130_fd_sc_hd__a21o_1 _1424_ (.A1(_0505_),
    .A2(_0716_),
    .B1(net66),
    .X(_0828_));
 sky130_fd_sc_hd__or2_2 _1425_ (.A(_0662_),
    .B(_0693_),
    .X(_0829_));
 sky130_fd_sc_hd__a22o_1 _1426_ (.A1(\cpu_inst.PC[0] ),
    .A2(_0820_),
    .B1(_0828_),
    .B2(net85),
    .X(_0830_));
 sky130_fd_sc_hd__a221o_1 _1427_ (.A1(\cpu_inst.C ),
    .A2(_0827_),
    .B1(_0829_),
    .B2(\cpu_inst.PC[8] ),
    .C1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__a221o_1 _1428_ (.A1(net4),
    .A2(net32),
    .B1(_0826_),
    .B2(_0831_),
    .C1(net16),
    .X(_0832_));
 sky130_fd_sc_hd__o22a_1 _1429_ (.A1(net99),
    .A2(net14),
    .B1(_0825_),
    .B2(_0832_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _1430_ (.A0(\cpu_inst.AXYS[3][1] ),
    .A1(\cpu_inst.AXYS[2][1] ),
    .S(net26),
    .X(_0833_));
 sky130_fd_sc_hd__and3_1 _1431_ (.A(\cpu_inst.AXYS[0][1] ),
    .B(net26),
    .C(_0810_),
    .X(_0834_));
 sky130_fd_sc_hd__a221o_2 _1432_ (.A1(\cpu_inst.AXYS[1][1] ),
    .A2(_0816_),
    .B1(_0833_),
    .B2(_0811_),
    .C1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__a22o_1 _1433_ (.A1(\cpu_inst.PC[1] ),
    .A2(_0820_),
    .B1(_0827_),
    .B2(\cpu_inst.Z ),
    .X(_0836_));
 sky130_fd_sc_hd__a221o_1 _1434_ (.A1(net84),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\cpu_inst.PC[9] ),
    .C1(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__a221o_1 _1435_ (.A1(net99),
    .A2(net32),
    .B1(_0826_),
    .B2(_0837_),
    .C1(net16),
    .X(_0838_));
 sky130_fd_sc_hd__a31o_1 _1436_ (.A1(net40),
    .A2(_0823_),
    .A3(_0835_),
    .B1(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o21a_1 _1437_ (.A1(net98),
    .A2(net14),
    .B1(_0839_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(\cpu_inst.AXYS[3][2] ),
    .A1(\cpu_inst.AXYS[2][2] ),
    .S(net27),
    .X(_0840_));
 sky130_fd_sc_hd__and3_1 _1439_ (.A(\cpu_inst.AXYS[0][2] ),
    .B(net26),
    .C(_0810_),
    .X(_0841_));
 sky130_fd_sc_hd__a221oi_4 _1440_ (.A1(\cpu_inst.AXYS[1][2] ),
    .A2(_0816_),
    .B1(_0840_),
    .B2(_0811_),
    .C1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__nor2_1 _1441_ (.A(_0824_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__a22o_1 _1442_ (.A1(\cpu_inst.I ),
    .A2(_0827_),
    .B1(_0828_),
    .B2(net83),
    .X(_0844_));
 sky130_fd_sc_hd__a221o_1 _1443_ (.A1(\cpu_inst.PC[2] ),
    .A2(_0820_),
    .B1(_0829_),
    .B2(\cpu_inst.PC[10] ),
    .C1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__o22a_1 _1444_ (.A1(net98),
    .A2(net69),
    .B1(net32),
    .B2(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__o22a_1 _1445_ (.A1(net97),
    .A2(net13),
    .B1(_0843_),
    .B2(_0846_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _1446_ (.A0(\cpu_inst.AXYS[3][3] ),
    .A1(\cpu_inst.AXYS[2][3] ),
    .S(net27),
    .X(_0847_));
 sky130_fd_sc_hd__o22a_1 _1447_ (.A1(\cpu_inst.AXYS[0][3] ),
    .A2(_0814_),
    .B1(_0817_),
    .B2(\cpu_inst.AXYS[1][3] ),
    .X(_0848_));
 sky130_fd_sc_hd__o21ai_2 _1448_ (.A1(_0810_),
    .A2(_0847_),
    .B1(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__nor2_1 _1449_ (.A(_0824_),
    .B(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__a22o_1 _1450_ (.A1(\cpu_inst.PC[3] ),
    .A2(_0820_),
    .B1(_0827_),
    .B2(\cpu_inst.D ),
    .X(_0851_));
 sky130_fd_sc_hd__a221o_1 _1451_ (.A1(net82),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\cpu_inst.PC[11] ),
    .C1(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__a221o_1 _1452_ (.A1(net97),
    .A2(net32),
    .B1(_0826_),
    .B2(_0852_),
    .C1(net16),
    .X(_0853_));
 sky130_fd_sc_hd__o22a_1 _1453_ (.A1(net96),
    .A2(net12),
    .B1(_0850_),
    .B2(_0853_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _1454_ (.A0(\cpu_inst.AXYS[3][4] ),
    .A1(\cpu_inst.AXYS[2][4] ),
    .S(net27),
    .X(_0854_));
 sky130_fd_sc_hd__o22a_1 _1455_ (.A1(\cpu_inst.AXYS[0][4] ),
    .A2(_0814_),
    .B1(_0817_),
    .B2(\cpu_inst.AXYS[1][4] ),
    .X(_0855_));
 sky130_fd_sc_hd__o21ai_2 _1456_ (.A1(_0810_),
    .A2(_0854_),
    .B1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__nor2_1 _1457_ (.A(_0824_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21a_1 _1458_ (.A1(net66),
    .A2(_0716_),
    .B1(net81),
    .X(_0858_));
 sky130_fd_sc_hd__nor3_1 _1459_ (.A(\cpu_inst.NMI_edge ),
    .B(net2),
    .C(_0686_),
    .Y(_0859_));
 sky130_fd_sc_hd__a221o_1 _1460_ (.A1(\cpu_inst.PC[4] ),
    .A2(_0820_),
    .B1(_0829_),
    .B2(\cpu_inst.PC[12] ),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a211o_1 _1461_ (.A1(\cpu_inst.php ),
    .A2(_0716_),
    .B1(_0858_),
    .C1(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__a221o_1 _1462_ (.A1(net96),
    .A2(net32),
    .B1(_0826_),
    .B2(_0861_),
    .C1(net16),
    .X(_0862_));
 sky130_fd_sc_hd__o22a_1 _1463_ (.A1(\cpu_inst.DI[4] ),
    .A2(net12),
    .B1(_0857_),
    .B2(_0862_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _1464_ (.A0(\cpu_inst.AXYS[3][5] ),
    .A1(\cpu_inst.AXYS[2][5] ),
    .S(net27),
    .X(_0863_));
 sky130_fd_sc_hd__o22a_1 _1465_ (.A1(\cpu_inst.AXYS[0][5] ),
    .A2(_0814_),
    .B1(_0817_),
    .B2(\cpu_inst.AXYS[1][5] ),
    .X(_0864_));
 sky130_fd_sc_hd__o21ai_1 _1466_ (.A1(_0810_),
    .A2(_0863_),
    .B1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__nor2_1 _1467_ (.A(_0824_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__o21a_1 _1468_ (.A1(net66),
    .A2(_0716_),
    .B1(net80),
    .X(_0867_));
 sky130_fd_sc_hd__a21o_1 _1469_ (.A1(\cpu_inst.PC[5] ),
    .A2(_0820_),
    .B1(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__a211o_1 _1470_ (.A1(\cpu_inst.PC[13] ),
    .A2(_0829_),
    .B1(_0827_),
    .C1(net32),
    .X(_0869_));
 sky130_fd_sc_hd__o22a_1 _1471_ (.A1(\cpu_inst.DI[4] ),
    .A2(net68),
    .B1(_0868_),
    .B2(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__o22a_1 _1472_ (.A1(\cpu_inst.DI[5] ),
    .A2(net12),
    .B1(_0866_),
    .B2(_0870_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1473_ (.A0(\cpu_inst.AXYS[3][6] ),
    .A1(\cpu_inst.AXYS[2][6] ),
    .S(net27),
    .X(_0871_));
 sky130_fd_sc_hd__o22a_1 _1474_ (.A1(\cpu_inst.AXYS[0][6] ),
    .A2(_0814_),
    .B1(_0817_),
    .B2(\cpu_inst.AXYS[1][6] ),
    .X(_0872_));
 sky130_fd_sc_hd__o21ai_2 _1475_ (.A1(_0810_),
    .A2(_0871_),
    .B1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_1 _1476_ (.A(_0824_),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__a22o_1 _1477_ (.A1(\cpu_inst.V ),
    .A2(_0827_),
    .B1(_0828_),
    .B2(net79),
    .X(_0875_));
 sky130_fd_sc_hd__a221o_1 _1478_ (.A1(\cpu_inst.PC[6] ),
    .A2(_0820_),
    .B1(_0829_),
    .B2(\cpu_inst.PC[14] ),
    .C1(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__o22a_1 _1479_ (.A1(\cpu_inst.DI[5] ),
    .A2(net69),
    .B1(net33),
    .B2(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__o22a_1 _1480_ (.A1(net95),
    .A2(net12),
    .B1(_0874_),
    .B2(_0877_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1481_ (.A0(\cpu_inst.AXYS[3][7] ),
    .A1(\cpu_inst.AXYS[2][7] ),
    .S(net27),
    .X(_0878_));
 sky130_fd_sc_hd__o22a_1 _1482_ (.A1(\cpu_inst.AXYS[0][7] ),
    .A2(_0814_),
    .B1(_0817_),
    .B2(\cpu_inst.AXYS[1][7] ),
    .X(_0879_));
 sky130_fd_sc_hd__o21ai_2 _1483_ (.A1(_0810_),
    .A2(_0878_),
    .B1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__nor2_1 _1484_ (.A(_0824_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__a22o_1 _1485_ (.A1(\cpu_inst.N ),
    .A2(_0827_),
    .B1(_0828_),
    .B2(net78),
    .X(_0882_));
 sky130_fd_sc_hd__a221o_1 _1486_ (.A1(\cpu_inst.PC[7] ),
    .A2(_0820_),
    .B1(_0829_),
    .B2(\cpu_inst.PC[15] ),
    .C1(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__o22a_1 _1487_ (.A1(net95),
    .A2(net68),
    .B1(net33),
    .B2(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__o22a_1 _1488_ (.A1(net94),
    .A2(net12),
    .B1(_0881_),
    .B2(_0884_),
    .X(_0021_));
 sky130_fd_sc_hd__nor3_4 _1489_ (.A(_0619_),
    .B(_0797_),
    .C(_0821_),
    .Y(_0885_));
 sky130_fd_sc_hd__or3_2 _1490_ (.A(_0619_),
    .B(_0797_),
    .C(_0821_),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_1 _1491_ (.A(_0819_),
    .B(_0885_),
    .Y(_0887_));
 sky130_fd_sc_hd__or2_1 _1492_ (.A(_0654_),
    .B(_0659_),
    .X(_0888_));
 sky130_fd_sc_hd__or4_1 _1493_ (.A(_0546_),
    .B(_0561_),
    .C(_0635_),
    .D(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__o21bai_4 _1494_ (.A1(\cpu_inst.state[5] ),
    .A2(_0538_),
    .B1_N(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__or3_1 _1495_ (.A(net52),
    .B(_0688_),
    .C(_0820_),
    .X(_0891_));
 sky130_fd_sc_hd__or3_2 _1496_ (.A(_0569_),
    .B(_0636_),
    .C(_0657_),
    .X(_0892_));
 sky130_fd_sc_hd__or4_1 _1497_ (.A(net53),
    .B(_0648_),
    .C(_0891_),
    .D(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__or2_1 _1498_ (.A(_0629_),
    .B(_0698_),
    .X(_0894_));
 sky130_fd_sc_hd__or3_1 _1499_ (.A(_0558_),
    .B(_0671_),
    .C(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__or3_4 _1500_ (.A(_0890_),
    .B(_0893_),
    .C(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__or3_4 _1501_ (.A(_0543_),
    .B(_0554_),
    .C(net60),
    .X(_0897_));
 sky130_fd_sc_hd__or3_4 _1502_ (.A(net66),
    .B(_0703_),
    .C(_0759_),
    .X(_0898_));
 sky130_fd_sc_hd__or2_4 _1503_ (.A(_0897_),
    .B(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__or2_4 _1504_ (.A(_0551_),
    .B(_0700_),
    .X(_0900_));
 sky130_fd_sc_hd__or2_1 _1505_ (.A(net56),
    .B(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__nor4_1 _1506_ (.A(_0886_),
    .B(_0896_),
    .C(_0899_),
    .D(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__or4_4 _1507_ (.A(_0886_),
    .B(_0896_),
    .C(_0899_),
    .D(_0901_),
    .X(_0903_));
 sky130_fd_sc_hd__and2_1 _1508_ (.A(net85),
    .B(net56),
    .X(_0904_));
 sky130_fd_sc_hd__a221o_1 _1509_ (.A1(\cpu_inst.ABL[0] ),
    .A2(_0899_),
    .B1(_0900_),
    .B2(net99),
    .C1(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__a211o_1 _1510_ (.A1(net85),
    .A2(_0896_),
    .B1(net7),
    .C1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__o22a_1 _1511_ (.A1(\cpu_inst.PC[0] ),
    .A2(_0903_),
    .B1(_0906_),
    .B2(_0887_),
    .X(_0907_));
 sky130_fd_sc_hd__or2_1 _1512_ (.A(net94),
    .B(net68),
    .X(_0908_));
 sky130_fd_sc_hd__o221a_1 _1513_ (.A1(net210),
    .A2(net12),
    .B1(_0907_),
    .B2(net33),
    .C1(_0908_),
    .X(_0022_));
 sky130_fd_sc_hd__a22o_1 _1514_ (.A1(\cpu_inst.ADD[1] ),
    .A2(net58),
    .B1(_0900_),
    .B2(net98),
    .X(_0909_));
 sky130_fd_sc_hd__a211o_1 _1515_ (.A1(\cpu_inst.ABL[1] ),
    .A2(_0899_),
    .B1(net7),
    .C1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _1516_ (.A1(_0835_),
    .A2(_0886_),
    .B1(_0896_),
    .B2(net84),
    .X(_0911_));
 sky130_fd_sc_hd__o22a_1 _1517_ (.A1(\cpu_inst.PC[1] ),
    .A2(_0903_),
    .B1(_0910_),
    .B2(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__or2_1 _1518_ (.A(net210),
    .B(net68),
    .X(_0913_));
 sky130_fd_sc_hd__o221a_1 _1519_ (.A1(net215),
    .A2(net12),
    .B1(_0912_),
    .B2(net33),
    .C1(_0913_),
    .X(_0023_));
 sky130_fd_sc_hd__a22o_1 _1520_ (.A1(net83),
    .A2(net57),
    .B1(_0900_),
    .B2(net97),
    .X(_0914_));
 sky130_fd_sc_hd__a211o_1 _1521_ (.A1(\cpu_inst.ABL[2] ),
    .A2(_0899_),
    .B1(net8),
    .C1(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a2bb2o_1 _1522_ (.A1_N(_0842_),
    .A2_N(_0885_),
    .B1(_0896_),
    .B2(net83),
    .X(_0916_));
 sky130_fd_sc_hd__o22a_1 _1523_ (.A1(\cpu_inst.PC[2] ),
    .A2(_0903_),
    .B1(_0915_),
    .B2(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__or2_1 _1524_ (.A(\spi_sram_master_inst.data[9] ),
    .B(net68),
    .X(_0918_));
 sky130_fd_sc_hd__o221a_1 _1525_ (.A1(net230),
    .A2(net12),
    .B1(_0917_),
    .B2(net34),
    .C1(_0918_),
    .X(_0024_));
 sky130_fd_sc_hd__a22o_1 _1526_ (.A1(net82),
    .A2(net57),
    .B1(_0900_),
    .B2(net96),
    .X(_0919_));
 sky130_fd_sc_hd__a211o_1 _1527_ (.A1(\cpu_inst.ABL[3] ),
    .A2(_0899_),
    .B1(net8),
    .C1(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__a2bb2o_1 _1528_ (.A1_N(_0849_),
    .A2_N(_0885_),
    .B1(_0896_),
    .B2(net82),
    .X(_0921_));
 sky130_fd_sc_hd__o22a_1 _1529_ (.A1(\cpu_inst.PC[3] ),
    .A2(_0903_),
    .B1(_0920_),
    .B2(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__or2_1 _1530_ (.A(net270),
    .B(net68),
    .X(_0923_));
 sky130_fd_sc_hd__o221a_1 _1531_ (.A1(net206),
    .A2(net12),
    .B1(_0922_),
    .B2(net34),
    .C1(_0923_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _1532_ (.A1(net81),
    .A2(net57),
    .B1(_0900_),
    .B2(\cpu_inst.DI[4] ),
    .X(_0924_));
 sky130_fd_sc_hd__a211o_1 _1533_ (.A1(\cpu_inst.ABL[4] ),
    .A2(_0899_),
    .B1(net8),
    .C1(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__a2bb2o_1 _1534_ (.A1_N(_0856_),
    .A2_N(_0885_),
    .B1(_0896_),
    .B2(net81),
    .X(_0926_));
 sky130_fd_sc_hd__o22a_1 _1535_ (.A1(\cpu_inst.PC[4] ),
    .A2(_0903_),
    .B1(_0925_),
    .B2(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__or2_1 _1536_ (.A(\spi_sram_master_inst.data[11] ),
    .B(net68),
    .X(_0928_));
 sky130_fd_sc_hd__o221a_1 _1537_ (.A1(net225),
    .A2(net13),
    .B1(_0927_),
    .B2(net34),
    .C1(_0928_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_1 _1538_ (.A1(net80),
    .A2(net57),
    .B1(_0900_),
    .B2(\cpu_inst.DI[5] ),
    .X(_0929_));
 sky130_fd_sc_hd__a211o_1 _1539_ (.A1(\cpu_inst.ABL[5] ),
    .A2(_0899_),
    .B1(net8),
    .C1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__a2bb2o_1 _1540_ (.A1_N(_0865_),
    .A2_N(_0885_),
    .B1(_0896_),
    .B2(net80),
    .X(_0931_));
 sky130_fd_sc_hd__o22a_1 _1541_ (.A1(\cpu_inst.PC[5] ),
    .A2(_0903_),
    .B1(_0930_),
    .B2(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__or2_1 _1542_ (.A(\spi_sram_master_inst.data[12] ),
    .B(net68),
    .X(_0933_));
 sky130_fd_sc_hd__o221a_1 _1543_ (.A1(net232),
    .A2(net13),
    .B1(_0932_),
    .B2(net34),
    .C1(_0933_),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_1 _1544_ (.A1(net79),
    .A2(net57),
    .B1(_0900_),
    .B2(net95),
    .X(_0934_));
 sky130_fd_sc_hd__a211o_1 _1545_ (.A1(\cpu_inst.ABL[6] ),
    .A2(_0899_),
    .B1(net8),
    .C1(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__a2bb2o_1 _1546_ (.A1_N(_0873_),
    .A2_N(_0885_),
    .B1(_0896_),
    .B2(net79),
    .X(_0936_));
 sky130_fd_sc_hd__o22a_1 _1547_ (.A1(\cpu_inst.PC[6] ),
    .A2(_0903_),
    .B1(_0935_),
    .B2(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__or2_1 _1548_ (.A(net272),
    .B(net68),
    .X(_0938_));
 sky130_fd_sc_hd__o221a_1 _1549_ (.A1(net222),
    .A2(net13),
    .B1(_0937_),
    .B2(net34),
    .C1(_0938_),
    .X(_0028_));
 sky130_fd_sc_hd__a22o_1 _1550_ (.A1(net78),
    .A2(net57),
    .B1(_0900_),
    .B2(net94),
    .X(_0939_));
 sky130_fd_sc_hd__a211o_1 _1551_ (.A1(\cpu_inst.ABL[7] ),
    .A2(_0899_),
    .B1(net8),
    .C1(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__a2bb2o_1 _1552_ (.A1_N(_0880_),
    .A2_N(_0885_),
    .B1(_0896_),
    .B2(\cpu_inst.ADD[7] ),
    .X(_0941_));
 sky130_fd_sc_hd__o22a_1 _1553_ (.A1(\cpu_inst.PC[7] ),
    .A2(_0903_),
    .B1(_0940_),
    .B2(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__or2_1 _1554_ (.A(net271),
    .B(net69),
    .X(_0943_));
 sky130_fd_sc_hd__o221a_1 _1555_ (.A1(net217),
    .A2(net12),
    .B1(_0942_),
    .B2(net33),
    .C1(_0943_),
    .X(_0029_));
 sky130_fd_sc_hd__a221o_1 _1556_ (.A1(net99),
    .A2(_0890_),
    .B1(_0897_),
    .B2(net85),
    .C1(_0886_),
    .X(_0944_));
 sky130_fd_sc_hd__o21a_1 _1557_ (.A1(net55),
    .A2(_0898_),
    .B1(\cpu_inst.ABH[0] ),
    .X(_0945_));
 sky130_fd_sc_hd__or4_1 _1558_ (.A(_0893_),
    .B(net7),
    .C(_0944_),
    .D(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__o21a_1 _1559_ (.A1(\cpu_inst.PC[8] ),
    .A2(_0903_),
    .B1(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__or2_1 _1560_ (.A(\spi_sram_master_inst.data[15] ),
    .B(net68),
    .X(_0948_));
 sky130_fd_sc_hd__o221a_1 _1561_ (.A1(net224),
    .A2(net14),
    .B1(_0947_),
    .B2(net35),
    .C1(_0948_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _1562_ (.A(\cpu_inst.ABH[1] ),
    .B(net55),
    .X(_0949_));
 sky130_fd_sc_hd__a221o_1 _1563_ (.A1(net84),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\cpu_inst.ABH[1] ),
    .C1(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__a221o_1 _1564_ (.A1(net98),
    .A2(_0890_),
    .B1(net7),
    .B2(\cpu_inst.PC[9] ),
    .C1(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__or2_1 _1565_ (.A(\spi_sram_master_inst.data[16] ),
    .B(net70),
    .X(_0952_));
 sky130_fd_sc_hd__o221a_1 _1566_ (.A1(net211),
    .A2(net14),
    .B1(_0951_),
    .B2(net32),
    .C1(_0952_),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _1567_ (.A(\cpu_inst.ABH[2] ),
    .B(net55),
    .X(_0953_));
 sky130_fd_sc_hd__a221o_1 _1568_ (.A1(net83),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\cpu_inst.ABH[2] ),
    .C1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__a221o_1 _1569_ (.A1(net97),
    .A2(_0890_),
    .B1(net7),
    .B2(\cpu_inst.PC[10] ),
    .C1(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__or2_1 _1570_ (.A(\spi_sram_master_inst.data[17] ),
    .B(net70),
    .X(_0956_));
 sky130_fd_sc_hd__o221a_1 _1571_ (.A1(net235),
    .A2(net14),
    .B1(_0955_),
    .B2(net32),
    .C1(_0956_),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _1572_ (.A(\cpu_inst.ABH[3] ),
    .B(net59),
    .X(_0957_));
 sky130_fd_sc_hd__a221o_1 _1573_ (.A1(net82),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\cpu_inst.ABH[3] ),
    .C1(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__a221o_1 _1574_ (.A1(net96),
    .A2(_0890_),
    .B1(net7),
    .B2(\cpu_inst.PC[11] ),
    .C1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__or2_1 _1575_ (.A(\spi_sram_master_inst.data[18] ),
    .B(net69),
    .X(_0960_));
 sky130_fd_sc_hd__o221a_1 _1576_ (.A1(net213),
    .A2(net13),
    .B1(_0959_),
    .B2(net35),
    .C1(_0960_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _1577_ (.A(\cpu_inst.ABH[4] ),
    .B(net56),
    .X(_0961_));
 sky130_fd_sc_hd__a221o_1 _1578_ (.A1(net81),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\cpu_inst.ABH[4] ),
    .C1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__a221o_1 _1579_ (.A1(\cpu_inst.DI[4] ),
    .A2(_0890_),
    .B1(net7),
    .B2(\cpu_inst.PC[12] ),
    .C1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__or2_1 _1580_ (.A(net213),
    .B(net69),
    .X(_0964_));
 sky130_fd_sc_hd__o221a_1 _1581_ (.A1(net216),
    .A2(net13),
    .B1(_0963_),
    .B2(net35),
    .C1(_0964_),
    .X(_0034_));
 sky130_fd_sc_hd__o21a_1 _1582_ (.A1(net56),
    .A2(_0898_),
    .B1(\cpu_inst.ABH[5] ),
    .X(_0965_));
 sky130_fd_sc_hd__a21o_1 _1583_ (.A1(net80),
    .A2(_0897_),
    .B1(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__a221o_1 _1584_ (.A1(\cpu_inst.DI[5] ),
    .A2(_0890_),
    .B1(net7),
    .B2(\cpu_inst.PC[13] ),
    .C1(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__or2_1 _1585_ (.A(net216),
    .B(net69),
    .X(_0968_));
 sky130_fd_sc_hd__o221a_1 _1586_ (.A1(net218),
    .A2(net13),
    .B1(_0967_),
    .B2(net35),
    .C1(_0968_),
    .X(_0035_));
 sky130_fd_sc_hd__o21a_1 _1587_ (.A1(net56),
    .A2(_0898_),
    .B1(\cpu_inst.ABH[6] ),
    .X(_0969_));
 sky130_fd_sc_hd__a21o_1 _1588_ (.A1(net79),
    .A2(_0897_),
    .B1(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__a221o_1 _1589_ (.A1(net95),
    .A2(_0890_),
    .B1(net7),
    .B2(\cpu_inst.PC[14] ),
    .C1(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__or2_1 _1590_ (.A(\spi_sram_master_inst.data[21] ),
    .B(net69),
    .X(_0972_));
 sky130_fd_sc_hd__o221a_1 _1591_ (.A1(net219),
    .A2(net13),
    .B1(_0971_),
    .B2(net34),
    .C1(_0972_),
    .X(_0036_));
 sky130_fd_sc_hd__o21a_1 _1592_ (.A1(net56),
    .A2(_0898_),
    .B1(\cpu_inst.ABH[7] ),
    .X(_0973_));
 sky130_fd_sc_hd__a21o_1 _1593_ (.A1(net78),
    .A2(_0897_),
    .B1(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__a221o_1 _1594_ (.A1(net94),
    .A2(_0890_),
    .B1(net7),
    .B2(\cpu_inst.PC[15] ),
    .C1(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__or2_1 _1595_ (.A(\spi_sram_master_inst.data[22] ),
    .B(net69),
    .X(_0976_));
 sky130_fd_sc_hd__o221a_1 _1596_ (.A1(\spi_sram_master_inst.data[23] ),
    .A2(net13),
    .B1(_0975_),
    .B2(net34),
    .C1(_0976_),
    .X(_0037_));
 sky130_fd_sc_hd__o31a_1 _1597_ (.A1(_0540_),
    .A2(_0543_),
    .A3(_0559_),
    .B1(\cpu_inst.store ),
    .X(_0977_));
 sky130_fd_sc_hd__nor2_1 _1598_ (.A(_0824_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__a221o_1 _1599_ (.A1(net166),
    .A2(net67),
    .B1(net15),
    .B2(net194),
    .C1(_0978_),
    .X(_0038_));
 sky130_fd_sc_hd__and3_1 _1600_ (.A(_0580_),
    .B(_0608_),
    .C(_0676_),
    .X(_0979_));
 sky130_fd_sc_hd__nand2_1 _1601_ (.A(net22),
    .B(_0594_),
    .Y(_0980_));
 sky130_fd_sc_hd__nor2_1 _1602_ (.A(_0615_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__and3_2 _1603_ (.A(net62),
    .B(_0594_),
    .C(_0613_),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_1 _1604_ (.A1(net250),
    .A2(net18),
    .B1(_0979_),
    .B2(_0981_),
    .X(_0039_));
 sky130_fd_sc_hd__or3_4 _1605_ (.A(_0568_),
    .B(_0703_),
    .C(_0759_),
    .X(_0983_));
 sky130_fd_sc_hd__nand2_4 _1606_ (.A(\cpu_inst.op[3] ),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__a221o_1 _1607_ (.A1(\cpu_inst.backwards ),
    .A2(net55),
    .B1(_0983_),
    .B2(\cpu_inst.op[2] ),
    .C1(_0822_),
    .X(_0985_));
 sky130_fd_sc_hd__inv_2 _1608_ (.A(net11),
    .Y(_0986_));
 sky130_fd_sc_hd__nor2_2 _1609_ (.A(_0984_),
    .B(net10),
    .Y(_0987_));
 sky130_fd_sc_hd__or2_2 _1610_ (.A(_0638_),
    .B(_0680_),
    .X(_0988_));
 sky130_fd_sc_hd__nor3_1 _1611_ (.A(_0565_),
    .B(_0759_),
    .C(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__or2_1 _1612_ (.A(_0619_),
    .B(_0688_),
    .X(_0990_));
 sky130_fd_sc_hd__nor3_1 _1613_ (.A(_0695_),
    .B(_0821_),
    .C(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__or3_1 _1614_ (.A(_0629_),
    .B(net53),
    .C(_0648_),
    .X(_0992_));
 sky130_fd_sc_hd__or4_1 _1615_ (.A(net55),
    .B(_0648_),
    .C(net52),
    .D(_0797_),
    .X(_0993_));
 sky130_fd_sc_hd__or2_4 _1616_ (.A(net61),
    .B(_0703_),
    .X(_0994_));
 sky130_fd_sc_hd__nor4_1 _1617_ (.A(_0665_),
    .B(_0992_),
    .C(_0993_),
    .D(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__and3_2 _1618_ (.A(_0989_),
    .B(_0991_),
    .C(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__a22o_1 _1619_ (.A1(\cpu_inst.PC[6] ),
    .A2(net61),
    .B1(_0996_),
    .B2(net95),
    .X(_0997_));
 sky130_fd_sc_hd__o21ai_1 _1620_ (.A1(net10),
    .A2(_0997_),
    .B1(_0984_),
    .Y(_0998_));
 sky130_fd_sc_hd__a21oi_1 _1621_ (.A1(net10),
    .A2(_0997_),
    .B1(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__and2_2 _1622_ (.A(\cpu_inst.shift_right ),
    .B(_0983_),
    .X(_1000_));
 sky130_fd_sc_hd__nand2_4 _1623_ (.A(\cpu_inst.shift_right ),
    .B(_0983_),
    .Y(_1001_));
 sky130_fd_sc_hd__and2b_1 _1624_ (.A_N(\cpu_inst.load_only ),
    .B(_0568_),
    .X(_1002_));
 sky130_fd_sc_hd__nor2_1 _1625_ (.A(_0802_),
    .B(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__and3_4 _1626_ (.A(_0885_),
    .B(_0989_),
    .C(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__inv_2 _1627_ (.A(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(_0873_),
    .B(_1004_),
    .Y(_1006_));
 sky130_fd_sc_hd__or2_4 _1629_ (.A(_0891_),
    .B(_0992_),
    .X(_1007_));
 sky130_fd_sc_hd__a221o_1 _1630_ (.A1(\cpu_inst.ABH[6] ),
    .A2(net57),
    .B1(_1007_),
    .B2(\cpu_inst.ADD[6] ),
    .C1(_1006_),
    .X(_1008_));
 sky130_fd_sc_hd__a21oi_1 _1631_ (.A1(net95),
    .A2(_0994_),
    .B1(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__nand2_1 _1632_ (.A(\cpu_inst.op[0] ),
    .B(_0983_),
    .Y(_1010_));
 sky130_fd_sc_hd__o31a_2 _1633_ (.A1(_0556_),
    .A2(net64),
    .A3(_0983_),
    .B1(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__and3_2 _1634_ (.A(\cpu_inst.op[1] ),
    .B(_0983_),
    .C(_1010_),
    .X(_1012_));
 sky130_fd_sc_hd__nor2_2 _1635_ (.A(\cpu_inst.op[1] ),
    .B(_1010_),
    .Y(_1013_));
 sky130_fd_sc_hd__or2_1 _1636_ (.A(\cpu_inst.op[1] ),
    .B(_1010_),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _1637_ (.A0(_1013_),
    .A1(_1012_),
    .S(_0997_),
    .X(_1015_));
 sky130_fd_sc_hd__nand2_1 _1638_ (.A(_0997_),
    .B(_1011_),
    .Y(_1016_));
 sky130_fd_sc_hd__mux2_1 _1639_ (.A0(_1015_),
    .A1(_1016_),
    .S(_1009_),
    .X(_1017_));
 sky130_fd_sc_hd__nor2_1 _1640_ (.A(_0880_),
    .B(_1004_),
    .Y(_1018_));
 sky130_fd_sc_hd__a22o_1 _1641_ (.A1(\cpu_inst.ABH[7] ),
    .A2(net56),
    .B1(_0994_),
    .B2(net94),
    .X(_1019_));
 sky130_fd_sc_hd__a211o_1 _1642_ (.A1(net78),
    .A2(_1007_),
    .B1(_1018_),
    .C1(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__nand2_1 _1643_ (.A(_1000_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__o21ai_1 _1644_ (.A1(_1000_),
    .A2(_1017_),
    .B1(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__o21a_1 _1645_ (.A1(_0987_),
    .A2(_0999_),
    .B1(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _1646_ (.A1(\cpu_inst.PC[5] ),
    .A2(net61),
    .B1(_0996_),
    .B2(\cpu_inst.DI[5] ),
    .X(_1024_));
 sky130_fd_sc_hd__o21ai_1 _1647_ (.A1(net10),
    .A2(_1024_),
    .B1(_0984_),
    .Y(_1025_));
 sky130_fd_sc_hd__a21oi_1 _1648_ (.A1(net10),
    .A2(_1024_),
    .B1(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_1 _1649_ (.A(_0865_),
    .B(_1004_),
    .Y(_1027_));
 sky130_fd_sc_hd__a22o_1 _1650_ (.A1(\cpu_inst.ABH[5] ),
    .A2(net58),
    .B1(_0994_),
    .B2(\cpu_inst.DI[5] ),
    .X(_1028_));
 sky130_fd_sc_hd__a211o_1 _1651_ (.A1(net80),
    .A2(_1007_),
    .B1(_1027_),
    .C1(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__a21o_1 _1652_ (.A1(_1011_),
    .A2(_1024_),
    .B1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__mux2_1 _1653_ (.A0(_1013_),
    .A1(_1012_),
    .S(_1024_),
    .X(_1031_));
 sky130_fd_sc_hd__nand2_1 _1654_ (.A(_1029_),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__nor2_1 _1655_ (.A(_1001_),
    .B(_1009_),
    .Y(_1033_));
 sky130_fd_sc_hd__a31o_1 _1656_ (.A1(_1001_),
    .A2(_1030_),
    .A3(_1032_),
    .B1(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__o21a_1 _1657_ (.A1(_0987_),
    .A2(_1026_),
    .B1(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__a22o_1 _1658_ (.A1(\cpu_inst.PC[4] ),
    .A2(net61),
    .B1(_0996_),
    .B2(\cpu_inst.DI[4] ),
    .X(_1036_));
 sky130_fd_sc_hd__o21ai_1 _1659_ (.A1(net10),
    .A2(_1036_),
    .B1(_0984_),
    .Y(_1037_));
 sky130_fd_sc_hd__a21oi_1 _1660_ (.A1(net10),
    .A2(_1036_),
    .B1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__a221o_1 _1661_ (.A1(\cpu_inst.DI[4] ),
    .A2(_0994_),
    .B1(_1007_),
    .B2(net81),
    .C1(_0961_),
    .X(_1039_));
 sky130_fd_sc_hd__o21ba_1 _1662_ (.A1(_0856_),
    .A2(_1004_),
    .B1_N(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _1663_ (.A0(_1013_),
    .A1(_1012_),
    .S(_1036_),
    .X(_1041_));
 sky130_fd_sc_hd__nor2_1 _1664_ (.A(_1040_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__a31o_1 _1665_ (.A1(_1011_),
    .A2(_1036_),
    .A3(_1040_),
    .B1(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _1666_ (.A0(_1029_),
    .A1(_1043_),
    .S(_1001_),
    .X(_1044_));
 sky130_fd_sc_hd__o21ai_1 _1667_ (.A1(_0987_),
    .A2(_1038_),
    .B1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a22o_1 _1668_ (.A1(\cpu_inst.PC[2] ),
    .A2(net61),
    .B1(_0996_),
    .B2(net97),
    .X(_1046_));
 sky130_fd_sc_hd__o21ai_1 _1669_ (.A1(net10),
    .A2(_1046_),
    .B1(_0984_),
    .Y(_1047_));
 sky130_fd_sc_hd__a21oi_1 _1670_ (.A1(net10),
    .A2(_1046_),
    .B1(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__nor2_1 _1671_ (.A(_0987_),
    .B(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__nor2_1 _1672_ (.A(_0842_),
    .B(_1004_),
    .Y(_1050_));
 sky130_fd_sc_hd__a21o_1 _1673_ (.A1(net83),
    .A2(_1007_),
    .B1(_0953_),
    .X(_1051_));
 sky130_fd_sc_hd__a211o_1 _1674_ (.A1(net97),
    .A2(_0994_),
    .B1(_1050_),
    .C1(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(_1013_),
    .A1(_1012_),
    .S(_1046_),
    .X(_1053_));
 sky130_fd_sc_hd__nand2_1 _1676_ (.A(_1011_),
    .B(_1046_),
    .Y(_1054_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(_1054_),
    .A1(_1053_),
    .S(_1052_),
    .X(_1055_));
 sky130_fd_sc_hd__a221o_1 _1678_ (.A1(net96),
    .A2(_0994_),
    .B1(_1007_),
    .B2(net82),
    .C1(_0957_),
    .X(_1056_));
 sky130_fd_sc_hd__o21ba_1 _1679_ (.A1(_0849_),
    .A2(_1004_),
    .B1_N(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(_1055_),
    .A1(_1057_),
    .S(_1000_),
    .X(_1058_));
 sky130_fd_sc_hd__a22o_1 _1681_ (.A1(\cpu_inst.PC[1] ),
    .A2(net61),
    .B1(_0996_),
    .B2(net98),
    .X(_1059_));
 sky130_fd_sc_hd__o21ai_1 _1682_ (.A1(net11),
    .A2(_1059_),
    .B1(_0984_),
    .Y(_1060_));
 sky130_fd_sc_hd__a21oi_1 _1683_ (.A1(net11),
    .A2(_1059_),
    .B1(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__nor2_1 _1684_ (.A(_0987_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a221o_1 _1685_ (.A1(net98),
    .A2(_0994_),
    .B1(_1007_),
    .B2(net84),
    .C1(_0949_),
    .X(_1063_));
 sky130_fd_sc_hd__a21oi_1 _1686_ (.A1(_0835_),
    .A2(_1005_),
    .B1(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__a21o_1 _1687_ (.A1(_0835_),
    .A2(_1005_),
    .B1(_1063_),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _1688_ (.A0(_1013_),
    .A1(_1012_),
    .S(_1059_),
    .X(_1066_));
 sky130_fd_sc_hd__a21oi_1 _1689_ (.A1(_1011_),
    .A2(_1059_),
    .B1(_1065_),
    .Y(_1067_));
 sky130_fd_sc_hd__a21o_1 _1690_ (.A1(_1065_),
    .A2(_1066_),
    .B1(_1000_),
    .X(_1068_));
 sky130_fd_sc_hd__o2bb2a_1 _1691_ (.A1_N(_1000_),
    .A2_N(_1052_),
    .B1(_1067_),
    .B2(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__a31o_1 _1692_ (.A1(_0813_),
    .A2(_0815_),
    .A3(_0818_),
    .B1(_1004_),
    .X(_1070_));
 sky130_fd_sc_hd__a22o_1 _1693_ (.A1(\cpu_inst.ABH[0] ),
    .A2(net59),
    .B1(_0994_),
    .B2(net99),
    .X(_1071_));
 sky130_fd_sc_hd__a21oi_1 _1694_ (.A1(net85),
    .A2(_1007_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__a22o_1 _1695_ (.A1(\cpu_inst.PC[0] ),
    .A2(net61),
    .B1(_0996_),
    .B2(net99),
    .X(_1073_));
 sky130_fd_sc_hd__nand2_1 _1696_ (.A(_1012_),
    .B(_1073_),
    .Y(_0186_));
 sky130_fd_sc_hd__a21oi_1 _1697_ (.A1(_1070_),
    .A2(_1072_),
    .B1(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__nand2_1 _1698_ (.A(_1011_),
    .B(_1073_),
    .Y(_0188_));
 sky130_fd_sc_hd__and3_1 _1699_ (.A(_1070_),
    .B(_1072_),
    .C(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__o21ai_1 _1700_ (.A1(_1014_),
    .A2(_1073_),
    .B1(_1001_),
    .Y(_0190_));
 sky130_fd_sc_hd__o32a_1 _1701_ (.A1(_0187_),
    .A2(_0189_),
    .A3(_0190_),
    .B1(_1064_),
    .B2(_1001_),
    .X(_0191_));
 sky130_fd_sc_hd__o21ai_1 _1702_ (.A1(net11),
    .A2(_1073_),
    .B1(_0984_),
    .Y(_0192_));
 sky130_fd_sc_hd__a21oi_1 _1703_ (.A1(net11),
    .A2(_1073_),
    .B1(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__nor2_1 _1704_ (.A(_0987_),
    .B(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__o211a_1 _1705_ (.A1(_0703_),
    .A2(_0759_),
    .B1(_0502_),
    .C1(\cpu_inst.inc ),
    .X(_0195_));
 sky130_fd_sc_hd__a21oi_1 _1706_ (.A1(\cpu_inst.C ),
    .A2(_1002_),
    .B1(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _1707_ (.A(\cpu_inst.shift ),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__or4_1 _1708_ (.A(_0638_),
    .B(_0690_),
    .C(_0700_),
    .D(_0990_),
    .X(_0198_));
 sky130_fd_sc_hd__a31o_1 _1709_ (.A1(\cpu_inst.compare ),
    .A2(_0502_),
    .A3(_0568_),
    .B1(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__o31a_1 _1710_ (.A1(_0546_),
    .A2(_0561_),
    .A3(net55),
    .B1(\cpu_inst.ALU.CO ),
    .X(_0200_));
 sky130_fd_sc_hd__a31o_1 _1711_ (.A1(\cpu_inst.C ),
    .A2(\cpu_inst.rotate ),
    .A3(_0983_),
    .B1(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__or4_2 _1712_ (.A(_0992_),
    .B(_0197_),
    .C(_0199_),
    .D(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__o211a_1 _1713_ (.A1(_0984_),
    .A2(_0986_),
    .B1(_1001_),
    .C1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _1714_ (.A0(_0194_),
    .A1(_0193_),
    .S(_0191_),
    .X(_0204_));
 sky130_fd_sc_hd__a2bb2o_1 _1715_ (.A1_N(_0191_),
    .A2_N(_0194_),
    .B1(_0203_),
    .B2(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1716_ (.A0(_1062_),
    .A1(_1061_),
    .S(_1069_),
    .X(_0206_));
 sky130_fd_sc_hd__a2bb2o_1 _1717_ (.A1_N(_1062_),
    .A2_N(_1069_),
    .B1(_0205_),
    .B2(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _1718_ (.A0(_1049_),
    .A1(_1048_),
    .S(_1058_),
    .X(_0208_));
 sky130_fd_sc_hd__o2bb2a_1 _1719_ (.A1_N(_0207_),
    .A2_N(_0208_),
    .B1(_1049_),
    .B2(_1058_),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _1720_ (.A1(\cpu_inst.PC[3] ),
    .A2(_0621_),
    .B1(_0996_),
    .B2(net96),
    .X(_0210_));
 sky130_fd_sc_hd__o21ai_1 _1721_ (.A1(net11),
    .A2(_0210_),
    .B1(_0984_),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_1 _1722_ (.A1(net10),
    .A2(_0210_),
    .B1(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _1723_ (.A(_0987_),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__mux2_1 _1724_ (.A0(_1013_),
    .A1(_1012_),
    .S(_0210_),
    .X(_0214_));
 sky130_fd_sc_hd__nand2_1 _1725_ (.A(_1011_),
    .B(_0210_),
    .Y(_0215_));
 sky130_fd_sc_hd__mux2_1 _1726_ (.A0(_0214_),
    .A1(_0215_),
    .S(_1057_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1727_ (.A0(_1040_),
    .A1(_0216_),
    .S(_1001_),
    .X(_0217_));
 sky130_fd_sc_hd__or2_1 _1728_ (.A(_0213_),
    .B(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(_0213_),
    .A1(_0212_),
    .S(_0217_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2b_1 _1730_ (.A_N(_0209_),
    .B(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__xor2_1 _1731_ (.A(_0209_),
    .B(_0219_),
    .X(_0221_));
 sky130_fd_sc_hd__xor2_1 _1732_ (.A(_0205_),
    .B(_0206_),
    .X(_0222_));
 sky130_fd_sc_hd__xor2_1 _1733_ (.A(_0207_),
    .B(_0208_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _1734_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _1735_ (.A(\cpu_inst.adc_bcd ),
    .B(_0568_),
    .Y(_0225_));
 sky130_fd_sc_hd__o311a_1 _1736_ (.A1(_0221_),
    .A2(_0224_),
    .A3(_0225_),
    .B1(_0220_),
    .C1(_0218_),
    .X(_0226_));
 sky130_fd_sc_hd__nor2_1 _1737_ (.A(_1038_),
    .B(_1044_),
    .Y(_0227_));
 sky130_fd_sc_hd__o21a_1 _1738_ (.A1(_1038_),
    .A2(_1044_),
    .B1(_1045_),
    .X(_0228_));
 sky130_fd_sc_hd__o21ai_1 _1739_ (.A1(_0226_),
    .A2(_0227_),
    .B1(_1045_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ba_1 _1740_ (.A1(_1026_),
    .A2(_1034_),
    .B1_N(_1035_),
    .X(_0230_));
 sky130_fd_sc_hd__a21o_1 _1741_ (.A1(_0229_),
    .A2(_0230_),
    .B1(_1035_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _1742_ (.A(_0999_),
    .B(_1022_),
    .X(_0232_));
 sky130_fd_sc_hd__and2b_1 _1743_ (.A_N(_1023_),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__a21oi_1 _1744_ (.A1(_0231_),
    .A2(_0232_),
    .B1(_1023_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _1745_ (.A(_1000_),
    .B(_0202_),
    .Y(_0235_));
 sky130_fd_sc_hd__a22o_1 _1746_ (.A1(\cpu_inst.PC[7] ),
    .A2(_0621_),
    .B1(_0996_),
    .B2(\cpu_inst.DI[7] ),
    .X(_0236_));
 sky130_fd_sc_hd__a21oi_1 _1747_ (.A1(_1011_),
    .A2(_0236_),
    .B1(_1020_),
    .Y(_0237_));
 sky130_fd_sc_hd__o21ai_1 _1748_ (.A1(_1014_),
    .A2(_0236_),
    .B1(_1001_),
    .Y(_0238_));
 sky130_fd_sc_hd__a311o_1 _1749_ (.A1(_1012_),
    .A2(_1020_),
    .A3(_0236_),
    .B1(_0237_),
    .C1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__o21ai_1 _1750_ (.A1(net11),
    .A2(_0236_),
    .B1(_0984_),
    .Y(_0240_));
 sky130_fd_sc_hd__a21o_1 _1751_ (.A1(net11),
    .A2(_0236_),
    .B1(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__and2b_1 _1752_ (.A_N(_0987_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__a21oi_1 _1753_ (.A1(_0235_),
    .A2(_0239_),
    .B1(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__and3_1 _1754_ (.A(_0235_),
    .B(_0239_),
    .C(_0241_),
    .X(_0244_));
 sky130_fd_sc_hd__nor2_1 _1755_ (.A(_0243_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__xnor2_1 _1756_ (.A(_0234_),
    .B(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__xnor2_1 _1757_ (.A(_0229_),
    .B(_0230_),
    .Y(_0247_));
 sky130_fd_sc_hd__xnor2_1 _1758_ (.A(_0231_),
    .B(_0233_),
    .Y(_0248_));
 sky130_fd_sc_hd__a21oi_1 _1759_ (.A1(_0247_),
    .A2(_0248_),
    .B1(_0225_),
    .Y(_0249_));
 sky130_fd_sc_hd__a21o_1 _1760_ (.A1(_0246_),
    .A2(_0249_),
    .B1(net33),
    .X(_0250_));
 sky130_fd_sc_hd__a21oi_1 _1761_ (.A1(_1070_),
    .A2(_1072_),
    .B1(_1001_),
    .Y(_0251_));
 sky130_fd_sc_hd__o21ba_1 _1762_ (.A1(_0234_),
    .A2(_0244_),
    .B1_N(_0243_),
    .X(_0252_));
 sky130_fd_sc_hd__xnor2_1 _1763_ (.A(_0251_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__o22a_1 _1764_ (.A1(\cpu_inst.ALU.CO ),
    .A2(net42),
    .B1(_0250_),
    .B2(_0253_),
    .X(_0040_));
 sky130_fd_sc_hd__xor2_1 _1765_ (.A(_0203_),
    .B(_0204_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _1766_ (.A0(net85),
    .A1(_0254_),
    .S(net41),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1767_ (.A0(\cpu_inst.ADD[1] ),
    .A1(_0222_),
    .S(net41),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1768_ (.A0(net83),
    .A1(_0223_),
    .S(net42),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_1 _1769_ (.A(net82),
    .B(net42),
    .Y(_0255_));
 sky130_fd_sc_hd__a21oi_1 _1770_ (.A1(net42),
    .A2(_0221_),
    .B1(_0255_),
    .Y(_0044_));
 sky130_fd_sc_hd__xnor2_1 _1771_ (.A(_0226_),
    .B(_0228_),
    .Y(_0256_));
 sky130_fd_sc_hd__mux2_1 _1772_ (.A0(net81),
    .A1(_0256_),
    .S(net42),
    .X(_0045_));
 sky130_fd_sc_hd__nor2_1 _1773_ (.A(net80),
    .B(net42),
    .Y(_0257_));
 sky130_fd_sc_hd__a21oi_1 _1774_ (.A1(net43),
    .A2(_0247_),
    .B1(_0257_),
    .Y(_0046_));
 sky130_fd_sc_hd__nand2_1 _1775_ (.A(net79),
    .B(net33),
    .Y(_0258_));
 sky130_fd_sc_hd__o21ai_1 _1776_ (.A1(net33),
    .A2(_0248_),
    .B1(_0258_),
    .Y(_0047_));
 sky130_fd_sc_hd__mux2_1 _1777_ (.A0(net78),
    .A1(_0246_),
    .S(net42),
    .X(_0048_));
 sky130_fd_sc_hd__nor2_1 _1778_ (.A(net252),
    .B(net42),
    .Y(_0259_));
 sky130_fd_sc_hd__a21oi_1 _1779_ (.A1(net42),
    .A2(_0226_),
    .B1(_0259_),
    .Y(_0049_));
 sky130_fd_sc_hd__mux2_1 _1780_ (.A0(net200),
    .A1(_1020_),
    .S(net42),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _1781_ (.A(_0668_),
    .B(_0821_),
    .X(_0260_));
 sky130_fd_sc_hd__o21ai_1 _1782_ (.A1(\cpu_inst.state[4] ),
    .A2(_0655_),
    .B1(_0667_),
    .Y(_0261_));
 sky130_fd_sc_hd__or4_1 _1783_ (.A(_0665_),
    .B(_0889_),
    .C(_0993_),
    .D(_0994_),
    .X(_0262_));
 sky130_fd_sc_hd__a211o_1 _1784_ (.A1(_0260_),
    .A2(_0261_),
    .B1(_0262_),
    .C1(_0705_),
    .X(_0263_));
 sky130_fd_sc_hd__or4_1 _1785_ (.A(_0630_),
    .B(_0634_),
    .C(_0682_),
    .D(_0695_),
    .X(_0264_));
 sky130_fd_sc_hd__or4_1 _1786_ (.A(_0657_),
    .B(_0660_),
    .C(_0670_),
    .D(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _1787_ (.A(_0537_),
    .B(net64),
    .X(_0266_));
 sky130_fd_sc_hd__or2_1 _1788_ (.A(net54),
    .B(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__or4_1 _1789_ (.A(net52),
    .B(_0688_),
    .C(_0265_),
    .D(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__or4_1 _1790_ (.A(_0565_),
    .B(_0638_),
    .C(_0700_),
    .D(_0759_),
    .X(_0269_));
 sky130_fd_sc_hd__or4_1 _1791_ (.A(_0568_),
    .B(net60),
    .C(_0894_),
    .D(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__or4_1 _1792_ (.A(_0539_),
    .B(_0543_),
    .C(_0569_),
    .D(_0619_),
    .X(_0271_));
 sky130_fd_sc_hd__or4_1 _1793_ (.A(_0535_),
    .B(_0555_),
    .C(_0270_),
    .D(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor3_1 _1794_ (.A(_0263_),
    .B(_0268_),
    .C(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__nor3_2 _1795_ (.A(_0777_),
    .B(_0988_),
    .C(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__mux2_1 _1796_ (.A0(\cpu_inst.ABH[0] ),
    .A1(_0947_),
    .S(net5),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1797_ (.A0(net248),
    .A1(_0951_),
    .S(net5),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1798_ (.A0(net251),
    .A1(_0955_),
    .S(net5),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1799_ (.A0(net239),
    .A1(_0959_),
    .S(net5),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1800_ (.A0(net246),
    .A1(_0963_),
    .S(net5),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1801_ (.A0(\cpu_inst.ABH[5] ),
    .A1(_0967_),
    .S(net5),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1802_ (.A0(\cpu_inst.ABH[6] ),
    .A1(_0971_),
    .S(net5),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1803_ (.A0(\cpu_inst.ABH[7] ),
    .A1(_0975_),
    .S(net5),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1804_ (.A0(net203),
    .A1(_0907_),
    .S(net5),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(net207),
    .A1(_0912_),
    .S(net5),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1806_ (.A0(net209),
    .A1(_0917_),
    .S(net6),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(net208),
    .A1(_0922_),
    .S(net6),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1808_ (.A0(net237),
    .A1(_0927_),
    .S(net6),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1809_ (.A0(net229),
    .A1(_0932_),
    .S(net6),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(net227),
    .A1(_0937_),
    .S(net6),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1811_ (.A0(net247),
    .A1(_0942_),
    .S(net6),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1812_ (.A0(net94),
    .A1(\cpu_inst.backwards ),
    .S(net32),
    .X(_0067_));
 sky130_fd_sc_hd__or3_1 _1813_ (.A(\cpu_inst.shift ),
    .B(\cpu_inst.adc_sbc ),
    .C(\cpu_inst.compare ),
    .X(_0275_));
 sky130_fd_sc_hd__or4_1 _1814_ (.A(net91),
    .B(\cpu_inst.clc ),
    .C(\cpu_inst.plp ),
    .D(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__a2bb2o_1 _1815_ (.A1_N(\cpu_inst.write_back ),
    .A2_N(_0573_),
    .B1(net66),
    .B2(\cpu_inst.shift ),
    .X(_0277_));
 sky130_fd_sc_hd__o22a_1 _1816_ (.A1(\cpu_inst.sec ),
    .A2(_0276_),
    .B1(_0277_),
    .B2(net53),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _1817_ (.A0(_0498_),
    .A1(net85),
    .S(\cpu_inst.plp ),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _1818_ (.A0(_0279_),
    .A1(\cpu_inst.ALU.CO ),
    .S(_0275_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(_0280_),
    .A1(net99),
    .S(net53),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _1820_ (.A0(\cpu_inst.C ),
    .A1(_0281_),
    .S(_0278_),
    .X(_0068_));
 sky130_fd_sc_hd__a2111o_1 _1821_ (.A1(\cpu_inst.load_reg ),
    .A2(_0817_),
    .B1(_0573_),
    .C1(\cpu_inst.compare ),
    .D1(\cpu_inst.plp ),
    .X(_0282_));
 sky130_fd_sc_hd__o21a_1 _1822_ (.A1(\cpu_inst.bit_ins ),
    .A2(_0282_),
    .B1(_0267_),
    .X(_0283_));
 sky130_fd_sc_hd__o21ba_1 _1823_ (.A1(\cpu_inst.plp ),
    .A2(net53),
    .B1_N(net66),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _1824_ (.A0(net84),
    .A1(\cpu_inst.DI[1] ),
    .S(net53),
    .X(_0285_));
 sky130_fd_sc_hd__or4_1 _1825_ (.A(net83),
    .B(net84),
    .C(net85),
    .D(net78),
    .X(_0286_));
 sky130_fd_sc_hd__or4_1 _1826_ (.A(net80),
    .B(net79),
    .C(net81),
    .D(net82),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_1 _1827_ (.A(_0286_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__mux2_1 _1828_ (.A0(_0288_),
    .A1(_0285_),
    .S(_0284_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(net204),
    .A1(_0289_),
    .S(_0283_),
    .X(_0069_));
 sky130_fd_sc_hd__a211o_1 _1830_ (.A1(\cpu_inst.bit_ins ),
    .A2(_0568_),
    .B1(net64),
    .C1(net53),
    .X(_0290_));
 sky130_fd_sc_hd__o21ai_1 _1831_ (.A1(net66),
    .A2(_0290_),
    .B1(_0282_),
    .Y(_0291_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(net94),
    .A1(net78),
    .S(_0266_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(_0292_),
    .A1(net238),
    .S(_0291_),
    .X(_0070_));
 sky130_fd_sc_hd__or4_1 _1834_ (.A(\cpu_inst.plp ),
    .B(\cpu_inst.cld ),
    .C(\cpu_inst.sed ),
    .D(_0573_),
    .X(_0293_));
 sky130_fd_sc_hd__o21a_1 _1835_ (.A1(net64),
    .A2(net53),
    .B1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1836_ (.A0(net82),
    .A1(_0504_),
    .S(_0499_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _1837_ (.A0(_0295_),
    .A1(net96),
    .S(net54),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(net254),
    .A1(_0296_),
    .S(_0294_),
    .X(_0071_));
 sky130_fd_sc_hd__o32a_1 _1839_ (.A1(\cpu_inst.cli ),
    .A2(\cpu_inst.sei ),
    .A3(_0545_),
    .B1(\cpu_inst.plp ),
    .B2(_0496_),
    .X(_0297_));
 sky130_fd_sc_hd__o31a_1 _1840_ (.A1(net64),
    .A2(net53),
    .A3(_0759_),
    .B1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _1841_ (.A0(net83),
    .A1(_0503_),
    .S(_0759_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _1842_ (.A0(_0299_),
    .A1(net97),
    .S(net53),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _1843_ (.A0(\cpu_inst.I ),
    .A1(_0300_),
    .S(_0298_),
    .X(_0301_));
 sky130_fd_sc_hd__or2_1 _1844_ (.A(_0682_),
    .B(_0301_),
    .X(_0072_));
 sky130_fd_sc_hd__o41a_1 _1845_ (.A1(\cpu_inst.adc_sbc ),
    .A2(\cpu_inst.plp ),
    .A3(\cpu_inst.clv ),
    .A4(_0573_),
    .B1(_0290_),
    .X(_0302_));
 sky130_fd_sc_hd__xnor2_1 _1846_ (.A(\cpu_inst.ALU.BI7 ),
    .B(\cpu_inst.ALU.AI7 ),
    .Y(_0303_));
 sky130_fd_sc_hd__xnor2_1 _1847_ (.A(\cpu_inst.ALU.CO ),
    .B(net78),
    .Y(_0304_));
 sky130_fd_sc_hd__a21oi_1 _1848_ (.A1(_0303_),
    .A2(_0304_),
    .B1(\cpu_inst.clv ),
    .Y(_0305_));
 sky130_fd_sc_hd__o2111a_1 _1849_ (.A1(_0303_),
    .A2(_0304_),
    .B1(_0305_),
    .C1(net64),
    .D1(_0499_),
    .X(_0306_));
 sky130_fd_sc_hd__and3_1 _1850_ (.A(\cpu_inst.plp ),
    .B(net79),
    .C(net64),
    .X(_0307_));
 sky130_fd_sc_hd__a211o_1 _1851_ (.A1(net95),
    .A2(_0573_),
    .B1(_0306_),
    .C1(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _1852_ (.A0(net243),
    .A1(_0308_),
    .S(_0302_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_4 _1853_ (.A(net100),
    .B(net39),
    .C(_0988_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _1854_ (.A0(net129),
    .A1(net99),
    .S(_0309_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1855_ (.A0(net165),
    .A1(net98),
    .S(_0309_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1856_ (.A0(net135),
    .A1(net97),
    .S(_0309_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1857_ (.A0(net163),
    .A1(net96),
    .S(_0309_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1858_ (.A0(net240),
    .A1(\cpu_inst.DI[4] ),
    .S(_0309_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1859_ (.A0(net155),
    .A1(\cpu_inst.DI[5] ),
    .S(_0309_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(net140),
    .A1(net95),
    .S(_0309_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1861_ (.A0(net176),
    .A1(net94),
    .S(_0309_),
    .X(_0081_));
 sky130_fd_sc_hd__a31o_1 _1862_ (.A1(net77),
    .A2(net1),
    .A3(net17),
    .B1(_0309_),
    .X(_0082_));
 sky130_fd_sc_hd__nor2_1 _1863_ (.A(_0585_),
    .B(_0745_),
    .Y(_0310_));
 sky130_fd_sc_hd__and2b_1 _1864_ (.A_N(_0594_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_1 _1865_ (.A(_0596_),
    .B(_0613_),
    .Y(_0312_));
 sky130_fd_sc_hd__or2_1 _1866_ (.A(_0596_),
    .B(_0613_),
    .X(_0313_));
 sky130_fd_sc_hd__nor2_2 _1867_ (.A(_0608_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__a211o_1 _1868_ (.A1(_0587_),
    .A2(_0314_),
    .B1(_0311_),
    .C1(_0676_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _1869_ (.A(_0609_),
    .B(_0982_),
    .Y(_0316_));
 sky130_fd_sc_hd__and3_1 _1870_ (.A(_0609_),
    .B(_0982_),
    .C(_0310_),
    .X(_0317_));
 sky130_fd_sc_hd__a31o_1 _1871_ (.A1(_0608_),
    .A2(_0749_),
    .A3(_0312_),
    .B1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__nand2_1 _1872_ (.A(_0578_),
    .B(_0312_),
    .Y(_0319_));
 sky130_fd_sc_hd__inv_2 _1873_ (.A(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__a31o_1 _1874_ (.A1(net50),
    .A2(_0310_),
    .A3(_0314_),
    .B1(net17),
    .X(_0321_));
 sky130_fd_sc_hd__a21oi_1 _1875_ (.A1(_0595_),
    .A2(_0608_),
    .B1(_0589_),
    .Y(_0322_));
 sky130_fd_sc_hd__nor2_1 _1876_ (.A(_0586_),
    .B(_0592_),
    .Y(_0323_));
 sky130_fd_sc_hd__a31o_1 _1877_ (.A1(net50),
    .A2(_0314_),
    .A3(_0323_),
    .B1(_0322_),
    .X(_0324_));
 sky130_fd_sc_hd__a211o_1 _1878_ (.A1(_0581_),
    .A2(_0315_),
    .B1(_0318_),
    .C1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__o22a_1 _1879_ (.A1(net260),
    .A2(net21),
    .B1(_0321_),
    .B2(_0325_),
    .X(_0083_));
 sky130_fd_sc_hd__a21bo_1 _1880_ (.A1(net170),
    .A2(_0573_),
    .B1_N(net1),
    .X(_0084_));
 sky130_fd_sc_hd__o2111a_1 _1881_ (.A1(_0577_),
    .A2(_0582_),
    .B1(_0604_),
    .C1(_0610_),
    .D1(_0312_),
    .X(_0326_));
 sky130_fd_sc_hd__a31o_1 _1882_ (.A1(_0595_),
    .A2(_0609_),
    .A3(_0676_),
    .B1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__or4_1 _1883_ (.A(_0585_),
    .B(net71),
    .C(_0745_),
    .D(_0319_),
    .X(_0328_));
 sky130_fd_sc_hd__or3b_1 _1884_ (.A(net19),
    .B(_0327_),
    .C_N(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__o22a_1 _1885_ (.A1(net137),
    .A2(net20),
    .B1(_0678_),
    .B2(_0329_),
    .X(_0085_));
 sky130_fd_sc_hd__a31o_1 _1886_ (.A1(_0577_),
    .A2(_0676_),
    .A3(_0982_),
    .B1(net17),
    .X(_0330_));
 sky130_fd_sc_hd__a211o_1 _1887_ (.A1(_0744_),
    .A2(_0314_),
    .B1(_0317_),
    .C1(_0327_),
    .X(_0331_));
 sky130_fd_sc_hd__o22a_1 _1888_ (.A1(net159),
    .A2(net22),
    .B1(_0330_),
    .B2(_0331_),
    .X(_0086_));
 sky130_fd_sc_hd__or3b_1 _1889_ (.A(_0313_),
    .B(net71),
    .C_N(_0582_),
    .X(_0332_));
 sky130_fd_sc_hd__o31a_1 _1890_ (.A1(_0585_),
    .A2(net71),
    .A3(_0319_),
    .B1(_0316_),
    .X(_0333_));
 sky130_fd_sc_hd__a21oi_1 _1891_ (.A1(_0332_),
    .A2(_0333_),
    .B1(_0605_),
    .Y(_0334_));
 sky130_fd_sc_hd__a31o_1 _1892_ (.A1(_0595_),
    .A2(_0609_),
    .A3(_0676_),
    .B1(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__o22a_1 _1893_ (.A1(net146),
    .A2(net20),
    .B1(_0321_),
    .B2(_0335_),
    .X(_0087_));
 sky130_fd_sc_hd__a31o_1 _1894_ (.A1(_0604_),
    .A2(_0719_),
    .A3(_0982_),
    .B1(net19),
    .X(_0336_));
 sky130_fd_sc_hd__a41o_1 _1895_ (.A1(_0594_),
    .A2(_0611_),
    .A3(_0615_),
    .A4(_0323_),
    .B1(_0318_),
    .X(_0337_));
 sky130_fd_sc_hd__o32a_1 _1896_ (.A1(_0335_),
    .A2(_0336_),
    .A3(_0337_),
    .B1(net20),
    .B2(net177),
    .X(_0088_));
 sky130_fd_sc_hd__nor2_1 _1897_ (.A(_0592_),
    .B(_0745_),
    .Y(_0338_));
 sky130_fd_sc_hd__a221o_1 _1898_ (.A1(net50),
    .A2(_0709_),
    .B1(_0320_),
    .B2(_0338_),
    .C1(_0591_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _1899_ (.A0(net172),
    .A1(_0339_),
    .S(net20),
    .X(_0089_));
 sky130_fd_sc_hd__o2111a_1 _1900_ (.A1(_0590_),
    .A2(_0323_),
    .B1(_0615_),
    .C1(_0611_),
    .D1(_0594_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1901_ (.A0(net223),
    .A1(_0340_),
    .S(net21),
    .X(_0090_));
 sky130_fd_sc_hd__and3_1 _1902_ (.A(net22),
    .B(_0313_),
    .C(_0338_),
    .X(_0341_));
 sky130_fd_sc_hd__a21o_1 _1903_ (.A1(net244),
    .A2(net17),
    .B1(_0341_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1904_ (.A0(net144),
    .A1(_0314_),
    .S(net22),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _1905_ (.A(_0607_),
    .B(_0982_),
    .C(_0338_),
    .X(_0342_));
 sky130_fd_sc_hd__o22a_1 _1906_ (.A1(net201),
    .A2(net22),
    .B1(_0330_),
    .B2(_0342_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _1907_ (.A(net18),
    .B(_0663_),
    .Y(_0343_));
 sky130_fd_sc_hd__and3_1 _1908_ (.A(_0590_),
    .B(net71),
    .C(_0613_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _1909_ (.A0(net261),
    .A1(_0344_),
    .S(_0343_),
    .X(_0094_));
 sky130_fd_sc_hd__or4b_1 _1910_ (.A(net19),
    .B(_0745_),
    .C(_0594_),
    .D_N(_0593_),
    .X(_0345_));
 sky130_fd_sc_hd__a21bo_1 _1911_ (.A1(net242),
    .A2(net19),
    .B1_N(_0345_),
    .X(_0095_));
 sky130_fd_sc_hd__and3_1 _1912_ (.A(\cpu_inst.D ),
    .B(_0596_),
    .C(_0344_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _1913_ (.A0(\cpu_inst.adc_bcd ),
    .A1(_0346_),
    .S(_0343_),
    .X(_0096_));
 sky130_fd_sc_hd__or3b_1 _1914_ (.A(net50),
    .B(_0605_),
    .C_N(_0585_),
    .X(_0347_));
 sky130_fd_sc_hd__o21ai_1 _1915_ (.A1(_0589_),
    .A2(_0607_),
    .B1(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__a22o_1 _1916_ (.A1(\cpu_inst.compare ),
    .A2(net18),
    .B1(_0981_),
    .B2(_0348_),
    .X(_0097_));
 sky130_fd_sc_hd__a22o_1 _1917_ (.A1(\cpu_inst.shift_right ),
    .A2(net17),
    .B1(_0618_),
    .B2(_0744_),
    .X(_0098_));
 sky130_fd_sc_hd__a32o_1 _1918_ (.A1(_0596_),
    .A2(net71),
    .A3(_0338_),
    .B1(_0311_),
    .B2(_0610_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _1919_ (.A0(net255),
    .A1(_0349_),
    .S(net22),
    .X(_0099_));
 sky130_fd_sc_hd__a211o_1 _1920_ (.A1(_0607_),
    .A2(_0614_),
    .B1(_0589_),
    .C1(_0595_),
    .X(_0350_));
 sky130_fd_sc_hd__and3_1 _1921_ (.A(_0596_),
    .B(_0615_),
    .C(_0744_),
    .X(_0351_));
 sky130_fd_sc_hd__or2_1 _1922_ (.A(net269),
    .B(net22),
    .X(_0352_));
 sky130_fd_sc_hd__o41a_1 _1923_ (.A1(net18),
    .A2(_0610_),
    .A3(_0350_),
    .A4(_0351_),
    .B1(_0352_),
    .X(_0100_));
 sky130_fd_sc_hd__o311a_1 _1924_ (.A1(_0592_),
    .A2(net71),
    .A3(_0745_),
    .B1(_0347_),
    .C1(_0589_),
    .X(_0353_));
 sky130_fd_sc_hd__nand2b_1 _1925_ (.A_N(_0353_),
    .B(_0982_),
    .Y(_0354_));
 sky130_fd_sc_hd__and4_1 _1926_ (.A(_0582_),
    .B(_0604_),
    .C(_0610_),
    .D(_0722_),
    .X(_0355_));
 sky130_fd_sc_hd__o211ai_1 _1927_ (.A1(_0677_),
    .A2(_0313_),
    .B1(_0350_),
    .C1(_0354_),
    .Y(_0356_));
 sky130_fd_sc_hd__a2111o_1 _1928_ (.A1(_0617_),
    .A2(_0744_),
    .B1(_0317_),
    .C1(_0355_),
    .D1(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__and3_1 _1929_ (.A(net23),
    .B(_0596_),
    .C(_0615_),
    .X(_0358_));
 sky130_fd_sc_hd__o2bb2a_1 _1930_ (.A1_N(_0357_),
    .A2_N(_0358_),
    .B1(\cpu_inst.op[1] ),
    .B2(net22),
    .X(_0101_));
 sky130_fd_sc_hd__or2_1 _1931_ (.A(net18),
    .B(_0357_),
    .X(_0359_));
 sky130_fd_sc_hd__o21a_1 _1932_ (.A1(net164),
    .A2(net22),
    .B1(_0359_),
    .X(_0102_));
 sky130_fd_sc_hd__o221a_1 _1933_ (.A1(\cpu_inst.op[3] ),
    .A2(net22),
    .B1(_0351_),
    .B2(_0359_),
    .C1(_0980_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1934_ (.A0(net236),
    .A1(_0355_),
    .S(net23),
    .X(_0104_));
 sky130_fd_sc_hd__and3_1 _1935_ (.A(_0580_),
    .B(_0676_),
    .C(_0314_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _1936_ (.A0(net249),
    .A1(_0360_),
    .S(net23),
    .X(_0105_));
 sky130_fd_sc_hd__and3_1 _1937_ (.A(_0580_),
    .B(net71),
    .C(_0676_),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _1938_ (.A1(net195),
    .A2(net17),
    .B1(_0618_),
    .B2(_0361_),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_1 _1939_ (.A1(net253),
    .A2(net17),
    .B1(_0618_),
    .B2(_0979_),
    .X(_0107_));
 sky130_fd_sc_hd__a22o_1 _1940_ (.A1(net174),
    .A2(net18),
    .B1(_0981_),
    .B2(_0361_),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_1 _1941_ (.A1(net190),
    .A2(net17),
    .B1(_0358_),
    .B2(_0361_),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _1942_ (.A1(net245),
    .A2(net17),
    .B1(_0979_),
    .B2(_0358_),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _1943_ (.A1(\cpu_inst.php ),
    .A2(net17),
    .B1(_0615_),
    .B2(_0679_),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _1944_ (.A1(\cpu_inst.plp ),
    .A2(net19),
    .B1(_0615_),
    .B2(_0727_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1945_ (.A0(net205),
    .A1(_0610_),
    .S(net39),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1946_ (.A0(net241),
    .A1(_0614_),
    .S(net39),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1947_ (.A0(net221),
    .A1(_0595_),
    .S(net39),
    .X(_0115_));
 sky130_fd_sc_hd__a211o_1 _1948_ (.A1(_0497_),
    .A2(_0531_),
    .B1(net61),
    .C1(_0682_),
    .X(_0362_));
 sky130_fd_sc_hd__a211o_1 _1949_ (.A1(net65),
    .A2(net62),
    .B1(_0757_),
    .C1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__or4_4 _1950_ (.A(_0674_),
    .B(_0705_),
    .C(_0888_),
    .D(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__or3_2 _1951_ (.A(_0535_),
    .B(_0635_),
    .C(_0888_),
    .X(_0365_));
 sky130_fd_sc_hd__or4_1 _1952_ (.A(net64),
    .B(net60),
    .C(net55),
    .D(net24),
    .X(_0366_));
 sky130_fd_sc_hd__a2bb2o_2 _1953_ (.A1_N(net52),
    .A2_N(_0366_),
    .B1(net65),
    .B2(net63),
    .X(_0367_));
 sky130_fd_sc_hd__or2_2 _1954_ (.A(net60),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__nor2_1 _1955_ (.A(_0573_),
    .B(net63),
    .Y(_0369_));
 sky130_fd_sc_hd__a221o_1 _1956_ (.A1(\cpu_inst.ADD[0] ),
    .A2(net24),
    .B1(net46),
    .B2(\cpu_inst.ABL[0] ),
    .C1(_0904_),
    .X(_0370_));
 sky130_fd_sc_hd__a21o_1 _1957_ (.A1(\cpu_inst.PC[0] ),
    .A2(_0368_),
    .B1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__xor2_1 _1958_ (.A(_0364_),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _1959_ (.A0(\cpu_inst.PC[0] ),
    .A1(_0372_),
    .S(net41),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_1 _1960_ (.A1(\cpu_inst.ADD[1] ),
    .A2(net58),
    .B1(net46),
    .B2(\cpu_inst.ABL[1] ),
    .X(_0373_));
 sky130_fd_sc_hd__a2bb2o_1 _1961_ (.A1_N(\cpu_inst.res ),
    .A2_N(_0686_),
    .B1(net24),
    .B2(net84),
    .X(_0374_));
 sky130_fd_sc_hd__a211o_1 _1962_ (.A1(\cpu_inst.PC[1] ),
    .A2(_0368_),
    .B1(_0373_),
    .C1(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__and3_1 _1963_ (.A(_0364_),
    .B(_0371_),
    .C(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__a21oi_1 _1964_ (.A1(_0364_),
    .A2(_0371_),
    .B1(_0375_),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_1 _1965_ (.A(_0376_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__mux2_1 _1966_ (.A0(\cpu_inst.PC[1] ),
    .A1(_0378_),
    .S(net41),
    .X(_0117_));
 sky130_fd_sc_hd__o21a_1 _1967_ (.A1(_0494_),
    .A2(\cpu_inst.res ),
    .B1(net52),
    .X(_0379_));
 sky130_fd_sc_hd__a221o_1 _1968_ (.A1(net83),
    .A2(net57),
    .B1(net47),
    .B2(\cpu_inst.ABL[2] ),
    .C1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__a221o_1 _1969_ (.A1(\cpu_inst.ADD[2] ),
    .A2(net25),
    .B1(_0368_),
    .B2(\cpu_inst.PC[2] ),
    .C1(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__xor2_1 _1970_ (.A(_0376_),
    .B(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _1971_ (.A0(net266),
    .A1(_0382_),
    .S(net43),
    .X(_0118_));
 sky130_fd_sc_hd__a221o_1 _1972_ (.A1(\cpu_inst.ADD[3] ),
    .A2(net57),
    .B1(net47),
    .B2(\cpu_inst.ABL[3] ),
    .C1(net51),
    .X(_0383_));
 sky130_fd_sc_hd__a221o_1 _1973_ (.A1(\cpu_inst.ADD[3] ),
    .A2(net25),
    .B1(_0368_),
    .B2(\cpu_inst.PC[3] ),
    .C1(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__a21oi_1 _1974_ (.A1(_0376_),
    .A2(_0381_),
    .B1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _1975_ (.A(_0376_),
    .B(_0381_),
    .C(_0384_),
    .X(_0386_));
 sky130_fd_sc_hd__nor2_1 _1976_ (.A(_0385_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__mux2_1 _1977_ (.A0(\cpu_inst.PC[3] ),
    .A1(_0387_),
    .S(net43),
    .X(_0119_));
 sky130_fd_sc_hd__a221o_1 _1978_ (.A1(net81),
    .A2(net57),
    .B1(net47),
    .B2(\cpu_inst.ABL[4] ),
    .C1(_0685_),
    .X(_0388_));
 sky130_fd_sc_hd__a221o_1 _1979_ (.A1(net81),
    .A2(net25),
    .B1(_0368_),
    .B2(\cpu_inst.PC[4] ),
    .C1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__xor2_1 _1980_ (.A(_0386_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _1981_ (.A0(net268),
    .A1(_0390_),
    .S(net43),
    .X(_0120_));
 sky130_fd_sc_hd__a221o_1 _1982_ (.A1(net80),
    .A2(net58),
    .B1(net47),
    .B2(\cpu_inst.ABL[5] ),
    .C1(_0685_),
    .X(_0391_));
 sky130_fd_sc_hd__a221o_1 _1983_ (.A1(net80),
    .A2(net25),
    .B1(_0368_),
    .B2(\cpu_inst.PC[5] ),
    .C1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__a21oi_1 _1984_ (.A1(_0386_),
    .A2(_0389_),
    .B1(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__and3_1 _1985_ (.A(_0386_),
    .B(_0389_),
    .C(_0392_),
    .X(_0394_));
 sky130_fd_sc_hd__nor2_1 _1986_ (.A(_0393_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__mux2_1 _1987_ (.A0(\cpu_inst.PC[5] ),
    .A1(_0395_),
    .S(net43),
    .X(_0121_));
 sky130_fd_sc_hd__a221o_1 _1988_ (.A1(net79),
    .A2(net58),
    .B1(net47),
    .B2(\cpu_inst.ABL[6] ),
    .C1(net51),
    .X(_0396_));
 sky130_fd_sc_hd__a221o_1 _1989_ (.A1(net79),
    .A2(net25),
    .B1(_0368_),
    .B2(\cpu_inst.PC[6] ),
    .C1(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__xor2_1 _1990_ (.A(_0394_),
    .B(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _1991_ (.A0(\cpu_inst.PC[6] ),
    .A1(_0398_),
    .S(net43),
    .X(_0122_));
 sky130_fd_sc_hd__a221o_1 _1992_ (.A1(\cpu_inst.ADD[7] ),
    .A2(net58),
    .B1(net47),
    .B2(\cpu_inst.ABL[7] ),
    .C1(net51),
    .X(_0399_));
 sky130_fd_sc_hd__a221o_1 _1993_ (.A1(\cpu_inst.ADD[7] ),
    .A2(net25),
    .B1(_0368_),
    .B2(\cpu_inst.PC[7] ),
    .C1(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__a21oi_1 _1994_ (.A1(_0394_),
    .A2(_0397_),
    .B1(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__and3_2 _1995_ (.A(_0394_),
    .B(_0397_),
    .C(_0400_),
    .X(_0402_));
 sky130_fd_sc_hd__nor2_1 _1996_ (.A(_0401_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__mux2_1 _1997_ (.A0(\cpu_inst.PC[7] ),
    .A1(_0403_),
    .S(net43),
    .X(_0123_));
 sky130_fd_sc_hd__a221o_1 _1998_ (.A1(net85),
    .A2(net60),
    .B1(net59),
    .B2(\cpu_inst.ABH[0] ),
    .C1(net52),
    .X(_0404_));
 sky130_fd_sc_hd__a221o_1 _1999_ (.A1(\cpu_inst.DI[0] ),
    .A2(net24),
    .B1(net46),
    .B2(\cpu_inst.ABH[0] ),
    .C1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__a21o_1 _2000_ (.A1(\cpu_inst.PC[8] ),
    .A2(_0367_),
    .B1(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__xor2_1 _2001_ (.A(_0402_),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _2002_ (.A0(net262),
    .A1(_0407_),
    .S(net40),
    .X(_0124_));
 sky130_fd_sc_hd__a211o_1 _2003_ (.A1(net84),
    .A2(net60),
    .B1(net52),
    .C1(_0949_),
    .X(_0408_));
 sky130_fd_sc_hd__a221o_1 _2004_ (.A1(net98),
    .A2(net24),
    .B1(net46),
    .B2(\cpu_inst.ABH[1] ),
    .C1(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__a21o_1 _2005_ (.A1(\cpu_inst.PC[9] ),
    .A2(_0367_),
    .B1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__a21oi_1 _2006_ (.A1(_0402_),
    .A2(_0406_),
    .B1(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__and3_1 _2007_ (.A(_0402_),
    .B(_0406_),
    .C(_0410_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _2008_ (.A(_0411_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__mux2_1 _2009_ (.A0(net258),
    .A1(_0413_),
    .S(net40),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _2010_ (.A1(net83),
    .A2(net60),
    .B1(net46),
    .B2(\cpu_inst.ABH[2] ),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _2011_ (.A1(net97),
    .A2(net24),
    .B1(_0367_),
    .B2(\cpu_inst.PC[10] ),
    .X(_0415_));
 sky130_fd_sc_hd__or4_1 _2012_ (.A(net51),
    .B(_0953_),
    .C(_0414_),
    .D(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__xor2_1 _2013_ (.A(_0412_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _2014_ (.A0(net267),
    .A1(_0417_),
    .S(net44),
    .X(_0126_));
 sky130_fd_sc_hd__a211o_1 _2015_ (.A1(net82),
    .A2(net60),
    .B1(net51),
    .C1(_0957_),
    .X(_0418_));
 sky130_fd_sc_hd__a221o_1 _2016_ (.A1(net96),
    .A2(net24),
    .B1(net46),
    .B2(\cpu_inst.ABH[3] ),
    .C1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__a21o_1 _2017_ (.A1(\cpu_inst.PC[11] ),
    .A2(_0367_),
    .B1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__a21oi_1 _2018_ (.A1(_0412_),
    .A2(_0416_),
    .B1(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__and3_1 _2019_ (.A(_0412_),
    .B(_0416_),
    .C(_0420_),
    .X(_0422_));
 sky130_fd_sc_hd__nor2_1 _2020_ (.A(_0421_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__mux2_1 _2021_ (.A0(net256),
    .A1(_0423_),
    .S(net44),
    .X(_0127_));
 sky130_fd_sc_hd__a211o_1 _2022_ (.A1(net81),
    .A2(_0642_),
    .B1(net51),
    .C1(_0961_),
    .X(_0424_));
 sky130_fd_sc_hd__a221o_1 _2023_ (.A1(\cpu_inst.DI[4] ),
    .A2(net24),
    .B1(net46),
    .B2(\cpu_inst.ABH[4] ),
    .C1(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__a21o_1 _2024_ (.A1(\cpu_inst.PC[12] ),
    .A2(_0367_),
    .B1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__xor2_1 _2025_ (.A(_0422_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _2026_ (.A0(net264),
    .A1(_0427_),
    .S(net41),
    .X(_0128_));
 sky130_fd_sc_hd__a221o_1 _2027_ (.A1(net80),
    .A2(_0642_),
    .B1(net56),
    .B2(\cpu_inst.ABH[5] ),
    .C1(net51),
    .X(_0428_));
 sky130_fd_sc_hd__a21o_1 _2028_ (.A1(\cpu_inst.ABH[5] ),
    .A2(net46),
    .B1(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__a221o_1 _2029_ (.A1(\cpu_inst.DI[5] ),
    .A2(net24),
    .B1(_0367_),
    .B2(\cpu_inst.PC[13] ),
    .C1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__a21oi_1 _2030_ (.A1(_0422_),
    .A2(_0426_),
    .B1(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__and3_1 _2031_ (.A(_0422_),
    .B(_0426_),
    .C(_0430_),
    .X(_0432_));
 sky130_fd_sc_hd__o21ai_1 _2032_ (.A1(_0431_),
    .A2(_0432_),
    .B1(net41),
    .Y(_0433_));
 sky130_fd_sc_hd__o21a_1 _2033_ (.A1(net259),
    .A2(net41),
    .B1(_0433_),
    .X(_0129_));
 sky130_fd_sc_hd__a221o_1 _2034_ (.A1(net79),
    .A2(_0642_),
    .B1(net56),
    .B2(\cpu_inst.ABH[6] ),
    .C1(net51),
    .X(_0434_));
 sky130_fd_sc_hd__a221o_1 _2035_ (.A1(\cpu_inst.DI[6] ),
    .A2(net25),
    .B1(net46),
    .B2(\cpu_inst.ABH[6] ),
    .C1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__a21o_1 _2036_ (.A1(\cpu_inst.PC[14] ),
    .A2(_0367_),
    .B1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__xor2_1 _2037_ (.A(_0432_),
    .B(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _2038_ (.A0(net265),
    .A1(_0437_),
    .S(net41),
    .X(_0130_));
 sky130_fd_sc_hd__a221o_1 _2039_ (.A1(net78),
    .A2(_0642_),
    .B1(net56),
    .B2(\cpu_inst.ABH[7] ),
    .C1(net51),
    .X(_0438_));
 sky130_fd_sc_hd__a221o_1 _2040_ (.A1(net94),
    .A2(net24),
    .B1(net46),
    .B2(\cpu_inst.ABH[7] ),
    .C1(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__a21o_1 _2041_ (.A1(\cpu_inst.PC[15] ),
    .A2(_0367_),
    .B1(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__and3_1 _2042_ (.A(_0432_),
    .B(_0436_),
    .C(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__a21oi_1 _2043_ (.A1(_0432_),
    .A2(_0436_),
    .B1(_0440_),
    .Y(_0442_));
 sky130_fd_sc_hd__o21ai_1 _2044_ (.A1(_0441_),
    .A2(_0442_),
    .B1(net41),
    .Y(_0443_));
 sky130_fd_sc_hd__o21a_1 _2045_ (.A1(net263),
    .A2(net41),
    .B1(_0443_),
    .X(_0131_));
 sky130_fd_sc_hd__or3b_1 _2046_ (.A(\cpu_inst.NMI_edge ),
    .B(net198),
    .C_N(net3),
    .X(_0444_));
 sky130_fd_sc_hd__o21ai_1 _2047_ (.A1(_0494_),
    .A2(_0682_),
    .B1(_0444_),
    .Y(_0132_));
 sky130_fd_sc_hd__a311o_1 _2048_ (.A1(_0499_),
    .A2(\cpu_inst.load_reg ),
    .A3(net64),
    .B1(_0682_),
    .C1(_0565_),
    .X(_0445_));
 sky130_fd_sc_hd__o31a_4 _2049_ (.A1(_0693_),
    .A2(_0892_),
    .A3(_0445_),
    .B1(net39),
    .X(_0446_));
 sky130_fd_sc_hd__nand3_4 _2050_ (.A(net26),
    .B(_0811_),
    .C(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__mux2_1 _2051_ (.A0(net99),
    .A1(net85),
    .S(_0694_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _2052_ (.A0(_0448_),
    .A1(net192),
    .S(_0447_),
    .X(_0133_));
 sky130_fd_sc_hd__and3_1 _2053_ (.A(\cpu_inst.adc_bcd ),
    .B(\cpu_inst.adj_bcd ),
    .C(\cpu_inst.ALU.HC ),
    .X(_0449_));
 sky130_fd_sc_hd__nand2b_1 _2054_ (.A_N(\cpu_inst.adc_bcd ),
    .B(\cpu_inst.adj_bcd ),
    .Y(_0450_));
 sky130_fd_sc_hd__nor2_1 _2055_ (.A(\cpu_inst.ALU.HC ),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__or3_1 _2056_ (.A(net84),
    .B(_0449_),
    .C(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__o21a_1 _2057_ (.A1(_0449_),
    .A2(_0451_),
    .B1(net84),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _2058_ (.A(_0693_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__a22o_1 _2059_ (.A1(net98),
    .A2(_0693_),
    .B1(_0452_),
    .B2(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _2060_ (.A0(_0455_),
    .A1(net156),
    .S(_0447_),
    .X(_0134_));
 sky130_fd_sc_hd__nand2_1 _2061_ (.A(\cpu_inst.ADD[2] ),
    .B(_0449_),
    .Y(_0456_));
 sky130_fd_sc_hd__or2_1 _2062_ (.A(\cpu_inst.ADD[2] ),
    .B(_0449_),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_1 _2063_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__xnor2_1 _2064_ (.A(_0453_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__mux2_1 _2065_ (.A0(\cpu_inst.DI[2] ),
    .A1(_0459_),
    .S(_0694_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(_0460_),
    .A1(net185),
    .S(_0447_),
    .X(_0135_));
 sky130_fd_sc_hd__a21bo_1 _2067_ (.A1(_0453_),
    .A2(_0457_),
    .B1_N(_0456_),
    .X(_0461_));
 sky130_fd_sc_hd__xnor2_1 _2068_ (.A(net82),
    .B(_0451_),
    .Y(_0462_));
 sky130_fd_sc_hd__xnor2_1 _2069_ (.A(_0461_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__mux2_1 _2070_ (.A0(\cpu_inst.DI[3] ),
    .A1(_0463_),
    .S(_0694_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _2071_ (.A0(_0464_),
    .A1(net187),
    .S(_0447_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(\cpu_inst.DI[4] ),
    .A1(\cpu_inst.ADD[4] ),
    .S(_0694_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _2073_ (.A0(_0465_),
    .A1(net173),
    .S(_0447_),
    .X(_0137_));
 sky130_fd_sc_hd__and3_1 _2074_ (.A(\cpu_inst.ALU.CO ),
    .B(\cpu_inst.adc_bcd ),
    .C(\cpu_inst.adj_bcd ),
    .X(_0466_));
 sky130_fd_sc_hd__nor2_1 _2075_ (.A(\cpu_inst.ALU.CO ),
    .B(_0450_),
    .Y(_0467_));
 sky130_fd_sc_hd__or3_1 _2076_ (.A(\cpu_inst.ADD[5] ),
    .B(_0466_),
    .C(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__o21a_1 _2077_ (.A1(_0466_),
    .A2(_0467_),
    .B1(\cpu_inst.ADD[5] ),
    .X(_0469_));
 sky130_fd_sc_hd__nor2_1 _2078_ (.A(_0693_),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__a22o_1 _2079_ (.A1(\cpu_inst.DI[5] ),
    .A2(_0693_),
    .B1(_0468_),
    .B2(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _2080_ (.A0(_0471_),
    .A1(net180),
    .S(_0447_),
    .X(_0138_));
 sky130_fd_sc_hd__nand2_1 _2081_ (.A(\cpu_inst.ADD[6] ),
    .B(_0466_),
    .Y(_0472_));
 sky130_fd_sc_hd__or2_1 _2082_ (.A(\cpu_inst.ADD[6] ),
    .B(_0466_),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _2083_ (.A(_0472_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__xnor2_1 _2084_ (.A(_0469_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__mux2_1 _2085_ (.A0(net95),
    .A1(_0475_),
    .S(_0694_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _2086_ (.A0(_0476_),
    .A1(net186),
    .S(_0447_),
    .X(_0139_));
 sky130_fd_sc_hd__a21bo_1 _2087_ (.A1(_0469_),
    .A2(_0473_),
    .B1_N(_0472_),
    .X(_0477_));
 sky130_fd_sc_hd__xnor2_1 _2088_ (.A(net78),
    .B(_0467_),
    .Y(_0478_));
 sky130_fd_sc_hd__xnor2_1 _2089_ (.A(_0477_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__mux2_1 _2090_ (.A0(\cpu_inst.DI[7] ),
    .A1(_0479_),
    .S(_0694_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _2091_ (.A0(_0480_),
    .A1(net179),
    .S(_0447_),
    .X(_0140_));
 sky130_fd_sc_hd__and3b_4 _2092_ (.A_N(net26),
    .B(_0811_),
    .C(_0446_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _2093_ (.A0(net184),
    .A1(_0448_),
    .S(_0481_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(net134),
    .A1(_0455_),
    .S(_0481_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2095_ (.A0(net133),
    .A1(_0460_),
    .S(_0481_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(net136),
    .A1(_0464_),
    .S(_0481_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2097_ (.A0(net131),
    .A1(_0465_),
    .S(_0481_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2098_ (.A0(net130),
    .A1(_0471_),
    .S(_0481_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2099_ (.A0(net132),
    .A1(_0476_),
    .S(_0481_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2100_ (.A0(net147),
    .A1(_0480_),
    .S(_0481_),
    .X(_0148_));
 sky130_fd_sc_hd__and3_4 _2101_ (.A(net26),
    .B(_0810_),
    .C(_0446_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _2102_ (.A0(net148),
    .A1(_0448_),
    .S(_0482_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2103_ (.A0(net143),
    .A1(_0455_),
    .S(_0482_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2104_ (.A0(net145),
    .A1(_0460_),
    .S(_0482_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2105_ (.A0(net168),
    .A1(_0464_),
    .S(_0482_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2106_ (.A0(net154),
    .A1(_0465_),
    .S(_0482_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(net161),
    .A1(_0471_),
    .S(_0482_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2108_ (.A0(net151),
    .A1(_0476_),
    .S(_0482_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(net183),
    .A1(_0480_),
    .S(_0482_),
    .X(_0156_));
 sky130_fd_sc_hd__a22o_1 _2110_ (.A1(\spi_sram_master_inst.data[23] ),
    .A2(net67),
    .B1(net16),
    .B2(net141),
    .X(_0157_));
 sky130_fd_sc_hd__a22o_1 _2111_ (.A1(net141),
    .A2(_0524_),
    .B1(net15),
    .B2(net189),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _2112_ (.A1(\spi_sram_master_inst.data[25] ),
    .A2(net67),
    .B1(net15),
    .B2(net149),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _2113_ (.A1(net149),
    .A2(net67),
    .B1(net16),
    .B2(net152),
    .X(_0160_));
 sky130_fd_sc_hd__a22o_1 _2114_ (.A1(net152),
    .A2(_0524_),
    .B1(net16),
    .B2(net160),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_1 _2115_ (.A1(net160),
    .A2(net67),
    .B1(net16),
    .B2(net171),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _2116_ (.A1(net171),
    .A2(_0524_),
    .B1(net15),
    .B2(net188),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_1 _2117_ (.A1(\spi_sram_master_inst.data[30] ),
    .A2(_0524_),
    .B1(net15),
    .B2(net166),
    .X(_0164_));
 sky130_fd_sc_hd__o22a_1 _2118_ (.A1(\spi_sram_master_inst.data[32] ),
    .A2(net70),
    .B1(net14),
    .B2(net126),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _2119_ (.A1(net126),
    .A2(net67),
    .B1(net15),
    .B2(net162),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _2120_ (.A1(\spi_sram_master_inst.data[34] ),
    .A2(net67),
    .B1(net15),
    .B2(net138),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _2121_ (.A1(net138),
    .A2(net67),
    .B1(net15),
    .B2(net153),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _2122_ (.A1(net153),
    .A2(net67),
    .B1(net15),
    .B2(net169),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _2123_ (.A1(\spi_sram_master_inst.data[37] ),
    .A2(net67),
    .B1(net15),
    .B2(net157),
    .X(_0170_));
 sky130_fd_sc_hd__o22a_1 _2124_ (.A1(\spi_sram_master_inst.data[38] ),
    .A2(net70),
    .B1(net14),
    .B2(net124),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_1 _2125_ (.A(\spi_sram_master_inst.counter_done ),
    .B(_0525_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_1 _2126_ (.A(_0506_),
    .B(_0514_),
    .Y(_0484_));
 sky130_fd_sc_hd__a211oi_1 _2127_ (.A1(\spi_sram_master_inst.state[1] ),
    .A2(\spi_sram_master_inst.counter_done ),
    .B1(_0507_),
    .C1(\spi_sram_master_inst.state[0] ),
    .Y(_0485_));
 sky130_fd_sc_hd__or3_1 _2128_ (.A(_0483_),
    .B(_0484_),
    .C(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__o21ai_1 _2129_ (.A1(_0484_),
    .A2(_0485_),
    .B1(_0483_),
    .Y(_0487_));
 sky130_fd_sc_hd__and3_1 _2130_ (.A(net100),
    .B(_0486_),
    .C(_0487_),
    .X(_0172_));
 sky130_fd_sc_hd__o311a_1 _2131_ (.A1(\spi_sram_master_inst.state[0] ),
    .A2(\spi_sram_master_inst.counter_done ),
    .A3(_0508_),
    .B1(_0510_),
    .C1(_0511_),
    .X(_0488_));
 sky130_fd_sc_hd__or3b_1 _2132_ (.A(_0483_),
    .B(_0484_),
    .C_N(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__o311a_1 _2133_ (.A1(\spi_sram_master_inst.state[1] ),
    .A2(\spi_sram_master_inst.counter_done ),
    .A3(_0525_),
    .B1(_0489_),
    .C1(net100),
    .X(_0173_));
 sky130_fd_sc_hd__a211o_1 _2134_ (.A1(\spi_sram_master_inst.state[2] ),
    .A2(_0483_),
    .B1(_0485_),
    .C1(_0520_),
    .X(_0490_));
 sky130_fd_sc_hd__and2_1 _2135_ (.A(net100),
    .B(_0490_),
    .X(_0174_));
 sky130_fd_sc_hd__and4_1 _2136_ (.A(\spi_sram_master_inst.state[1] ),
    .B(\spi_sram_master_inst.counter_done ),
    .C(net100),
    .D(_0506_),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _2137_ (.A(net33),
    .B(_0242_),
    .X(_0491_));
 sky130_fd_sc_hd__a2bb2o_1 _2138_ (.A1_N(_0244_),
    .A2_N(_0491_),
    .B1(net202),
    .B2(net33),
    .X(_0176_));
 sky130_fd_sc_hd__nand2_4 _2139_ (.A(_0816_),
    .B(_0446_),
    .Y(_0492_));
 sky130_fd_sc_hd__mux2_1 _2140_ (.A0(_0448_),
    .A1(net228),
    .S(_0492_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2141_ (.A0(_0455_),
    .A1(net182),
    .S(_0492_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2142_ (.A0(_0460_),
    .A1(net257),
    .S(_0492_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2143_ (.A0(_0464_),
    .A1(net175),
    .S(_0492_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2144_ (.A0(_0465_),
    .A1(net178),
    .S(_0492_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2145_ (.A0(_0471_),
    .A1(net181),
    .S(_0492_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2146_ (.A0(_0476_),
    .A1(net193),
    .S(_0492_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2147_ (.A0(_0480_),
    .A1(net191),
    .S(_0492_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _2149_ (.CLK(clknet_4_5_0_clk),
    .D(_0012_),
    .Q(\spi_sram_master_inst.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2150_ (.CLK(clknet_4_5_0_clk),
    .D(_0013_),
    .Q(\spi_sram_master_inst.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2151_ (.CLK(clknet_4_5_0_clk),
    .D(_0001_),
    .Q(\spi_sram_master_inst.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2152_ (.CLK(clknet_4_5_0_clk),
    .D(_0002_),
    .Q(\spi_sram_master_inst.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2153_ (.CLK(clknet_4_5_0_clk),
    .D(_0003_),
    .Q(\spi_sram_master_inst.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2154_ (.CLK(clknet_4_6_0_clk),
    .D(_0014_),
    .Q(\cpu_inst.DI[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2155_ (.CLK(clknet_4_3_0_clk),
    .D(_0015_),
    .Q(\cpu_inst.DI[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2156_ (.CLK(clknet_4_12_0_clk),
    .D(_0016_),
    .Q(\cpu_inst.DI[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2157_ (.CLK(clknet_4_14_0_clk),
    .D(_0017_),
    .Q(\cpu_inst.DI[3] ));
 sky130_fd_sc_hd__dfxtp_4 _2158_ (.CLK(clknet_4_14_0_clk),
    .D(_0018_),
    .Q(\cpu_inst.DI[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2159_ (.CLK(clknet_4_14_0_clk),
    .D(_0019_),
    .Q(\cpu_inst.DI[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2160_ (.CLK(clknet_4_14_0_clk),
    .D(_0020_),
    .Q(\cpu_inst.DI[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2161_ (.CLK(clknet_4_14_0_clk),
    .D(_0021_),
    .Q(\cpu_inst.DI[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2162_ (.CLK(clknet_4_15_0_clk),
    .D(_0022_),
    .Q(\spi_sram_master_inst.data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2163_ (.CLK(clknet_4_15_0_clk),
    .D(_0023_),
    .Q(\spi_sram_master_inst.data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2164_ (.CLK(clknet_4_15_0_clk),
    .D(net231),
    .Q(\spi_sram_master_inst.data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2165_ (.CLK(clknet_4_15_0_clk),
    .D(_0025_),
    .Q(\spi_sram_master_inst.data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2166_ (.CLK(clknet_4_15_0_clk),
    .D(net226),
    .Q(\spi_sram_master_inst.data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2167_ (.CLK(clknet_4_15_0_clk),
    .D(net233),
    .Q(\spi_sram_master_inst.data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2168_ (.CLK(clknet_4_15_0_clk),
    .D(_0028_),
    .Q(\spi_sram_master_inst.data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2169_ (.CLK(clknet_4_15_0_clk),
    .D(_0029_),
    .Q(\spi_sram_master_inst.data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2170_ (.CLK(clknet_4_6_0_clk),
    .D(_0030_),
    .Q(\spi_sram_master_inst.data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2171_ (.CLK(clknet_4_13_0_clk),
    .D(net212),
    .Q(\spi_sram_master_inst.data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2172_ (.CLK(clknet_4_13_0_clk),
    .D(_0032_),
    .Q(\spi_sram_master_inst.data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2173_ (.CLK(clknet_4_13_0_clk),
    .D(net214),
    .Q(\spi_sram_master_inst.data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2174_ (.CLK(clknet_4_13_0_clk),
    .D(_0034_),
    .Q(\spi_sram_master_inst.data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2175_ (.CLK(clknet_4_13_0_clk),
    .D(_0035_),
    .Q(\spi_sram_master_inst.data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2176_ (.CLK(clknet_4_13_0_clk),
    .D(net220),
    .Q(\spi_sram_master_inst.data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2177_ (.CLK(clknet_4_15_0_clk),
    .D(_0037_),
    .Q(\spi_sram_master_inst.data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2178_ (.CLK(clknet_4_7_0_clk),
    .D(_0038_),
    .Q(\spi_sram_master_inst.data[32] ));
 sky130_fd_sc_hd__dfrtp_1 _2179_ (.CLK(clknet_4_4_0_clk),
    .D(_0004_),
    .RESET_B(net100),
    .Q(\cpu_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2180_ (.CLK(clknet_4_1_0_clk),
    .D(_0005_),
    .RESET_B(net100),
    .Q(\cpu_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2181_ (.CLK(clknet_4_4_0_clk),
    .D(_0006_),
    .RESET_B(net100),
    .Q(\cpu_inst.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _2182_ (.CLK(clknet_4_4_0_clk),
    .D(_0007_),
    .SET_B(net100),
    .Q(\cpu_inst.state[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2183_ (.CLK(clknet_4_4_0_clk),
    .D(_0008_),
    .RESET_B(net100),
    .Q(\cpu_inst.state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2184_ (.CLK(clknet_4_4_0_clk),
    .D(_0009_),
    .RESET_B(net1),
    .Q(\cpu_inst.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2185_ (.CLK(clknet_4_2_0_clk),
    .D(_0039_),
    .Q(\cpu_inst.cld ));
 sky130_fd_sc_hd__dfxtp_4 _2186_ (.CLK(clknet_4_11_0_clk),
    .D(_0040_),
    .Q(\cpu_inst.ALU.CO ));
 sky130_fd_sc_hd__dfxtp_1 _2187_ (.CLK(clknet_4_9_0_clk),
    .D(_0041_),
    .Q(\cpu_inst.ADD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2188_ (.CLK(clknet_4_11_0_clk),
    .D(_0042_),
    .Q(\cpu_inst.ADD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2189_ (.CLK(clknet_4_11_0_clk),
    .D(_0043_),
    .Q(\cpu_inst.ADD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2190_ (.CLK(clknet_4_11_0_clk),
    .D(_0044_),
    .Q(\cpu_inst.ADD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2191_ (.CLK(clknet_4_11_0_clk),
    .D(_0045_),
    .Q(\cpu_inst.ADD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2192_ (.CLK(clknet_4_11_0_clk),
    .D(_0046_),
    .Q(\cpu_inst.ADD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2193_ (.CLK(clknet_4_11_0_clk),
    .D(_0047_),
    .Q(\cpu_inst.ADD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2194_ (.CLK(clknet_4_11_0_clk),
    .D(_0048_),
    .Q(\cpu_inst.ADD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2195_ (.CLK(clknet_4_11_0_clk),
    .D(_0049_),
    .Q(\cpu_inst.ALU.HC ));
 sky130_fd_sc_hd__dfxtp_1 _2196_ (.CLK(clknet_4_11_0_clk),
    .D(_0050_),
    .Q(\cpu_inst.ALU.AI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2197_ (.CLK(clknet_4_6_0_clk),
    .D(_0051_),
    .Q(\cpu_inst.ABH[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2198_ (.CLK(clknet_4_6_0_clk),
    .D(_0052_),
    .Q(\cpu_inst.ABH[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2199_ (.CLK(clknet_4_13_0_clk),
    .D(_0053_),
    .Q(\cpu_inst.ABH[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2200_ (.CLK(clknet_4_12_0_clk),
    .D(_0054_),
    .Q(\cpu_inst.ABH[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2201_ (.CLK(clknet_4_12_0_clk),
    .D(_0055_),
    .Q(\cpu_inst.ABH[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2202_ (.CLK(clknet_4_12_0_clk),
    .D(_0056_),
    .Q(\cpu_inst.ABH[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2203_ (.CLK(clknet_4_15_0_clk),
    .D(_0057_),
    .Q(\cpu_inst.ABH[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2204_ (.CLK(clknet_4_13_0_clk),
    .D(_0058_),
    .Q(\cpu_inst.ABH[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2205_ (.CLK(clknet_4_12_0_clk),
    .D(_0059_),
    .Q(\cpu_inst.ABL[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2206_ (.CLK(clknet_4_12_0_clk),
    .D(_0060_),
    .Q(\cpu_inst.ABL[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2207_ (.CLK(clknet_4_14_0_clk),
    .D(_0061_),
    .Q(\cpu_inst.ABL[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2208_ (.CLK(clknet_4_14_0_clk),
    .D(_0062_),
    .Q(\cpu_inst.ABL[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2209_ (.CLK(clknet_4_15_0_clk),
    .D(_0063_),
    .Q(\cpu_inst.ABL[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2210_ (.CLK(clknet_4_15_0_clk),
    .D(_0064_),
    .Q(\cpu_inst.ABL[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2211_ (.CLK(clknet_4_14_0_clk),
    .D(_0065_),
    .Q(\cpu_inst.ABL[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2212_ (.CLK(clknet_4_15_0_clk),
    .D(_0066_),
    .Q(\cpu_inst.ABL[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2213_ (.CLK(clknet_4_3_0_clk),
    .D(_0067_),
    .Q(\cpu_inst.backwards ));
 sky130_fd_sc_hd__dfxtp_1 _2214_ (.CLK(clknet_4_11_0_clk),
    .D(_0000_),
    .Q(\cpu_inst.adj_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2215_ (.CLK(clknet_4_3_0_clk),
    .D(_0068_),
    .Q(\cpu_inst.C ));
 sky130_fd_sc_hd__dfxtp_1 _2216_ (.CLK(clknet_4_9_0_clk),
    .D(_0069_),
    .Q(\cpu_inst.Z ));
 sky130_fd_sc_hd__dfxtp_1 _2217_ (.CLK(clknet_4_9_0_clk),
    .D(_0070_),
    .Q(\cpu_inst.N ));
 sky130_fd_sc_hd__dfxtp_1 _2218_ (.CLK(clknet_4_9_0_clk),
    .D(_0071_),
    .Q(\cpu_inst.D ));
 sky130_fd_sc_hd__dfxtp_1 _2219_ (.CLK(clknet_4_3_0_clk),
    .D(_0072_),
    .Q(\cpu_inst.I ));
 sky130_fd_sc_hd__dfxtp_1 _2220_ (.CLK(clknet_4_9_0_clk),
    .D(_0073_),
    .Q(\cpu_inst.V ));
 sky130_fd_sc_hd__dfxtp_1 _2221_ (.CLK(clknet_4_2_0_clk),
    .D(_0074_),
    .Q(\cpu_inst.IRHOLD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2222_ (.CLK(clknet_4_8_0_clk),
    .D(_0075_),
    .Q(\cpu_inst.IRHOLD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2223_ (.CLK(clknet_4_2_0_clk),
    .D(_0076_),
    .Q(\cpu_inst.IRHOLD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2224_ (.CLK(clknet_4_8_0_clk),
    .D(_0077_),
    .Q(\cpu_inst.IRHOLD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2225_ (.CLK(clknet_4_2_0_clk),
    .D(_0078_),
    .Q(\cpu_inst.IRHOLD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2226_ (.CLK(clknet_4_8_0_clk),
    .D(_0079_),
    .Q(\cpu_inst.IRHOLD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2227_ (.CLK(clknet_4_9_0_clk),
    .D(_0080_),
    .Q(\cpu_inst.IRHOLD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2228_ (.CLK(clknet_4_8_0_clk),
    .D(_0081_),
    .Q(\cpu_inst.IRHOLD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2229_ (.CLK(clknet_4_8_0_clk),
    .D(_0082_),
    .Q(\cpu_inst.IRHOLD_valid ));
 sky130_fd_sc_hd__dfxtp_1 _2230_ (.CLK(clknet_4_0_0_clk),
    .D(_0083_),
    .Q(\cpu_inst.load_reg ));
 sky130_fd_sc_hd__dfxtp_1 _2231_ (.CLK(clknet_4_6_0_clk),
    .D(_0084_),
    .Q(\cpu_inst.res ));
 sky130_fd_sc_hd__dfxtp_1 _2232_ (.CLK(clknet_4_0_0_clk),
    .D(_0085_),
    .Q(\cpu_inst.dst_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2233_ (.CLK(clknet_4_2_0_clk),
    .D(_0086_),
    .Q(\cpu_inst.dst_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2234_ (.CLK(clknet_4_0_0_clk),
    .D(_0087_),
    .Q(\cpu_inst.src_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2235_ (.CLK(clknet_4_0_0_clk),
    .D(_0088_),
    .Q(\cpu_inst.src_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2236_ (.CLK(clknet_4_0_0_clk),
    .D(_0089_),
    .Q(\cpu_inst.index_y ));
 sky130_fd_sc_hd__dfxtp_1 _2237_ (.CLK(clknet_4_1_0_clk),
    .D(_0090_),
    .Q(\cpu_inst.store ));
 sky130_fd_sc_hd__dfxtp_1 _2238_ (.CLK(clknet_4_0_0_clk),
    .D(_0091_),
    .Q(\cpu_inst.write_back ));
 sky130_fd_sc_hd__dfxtp_1 _2239_ (.CLK(clknet_4_2_0_clk),
    .D(_0092_),
    .Q(\cpu_inst.load_only ));
 sky130_fd_sc_hd__dfxtp_1 _2240_ (.CLK(clknet_4_2_0_clk),
    .D(_0093_),
    .Q(\cpu_inst.inc ));
 sky130_fd_sc_hd__dfxtp_1 _2241_ (.CLK(clknet_4_9_0_clk),
    .D(_0094_),
    .Q(\cpu_inst.adc_sbc ));
 sky130_fd_sc_hd__dfxtp_1 _2242_ (.CLK(clknet_4_0_0_clk),
    .D(_0095_),
    .Q(\cpu_inst.shift ));
 sky130_fd_sc_hd__dfxtp_1 _2243_ (.CLK(clknet_4_9_0_clk),
    .D(_0096_),
    .Q(\cpu_inst.adc_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2244_ (.CLK(clknet_4_2_0_clk),
    .D(_0097_),
    .Q(\cpu_inst.compare ));
 sky130_fd_sc_hd__dfxtp_1 _2245_ (.CLK(clknet_4_1_0_clk),
    .D(_0098_),
    .Q(\cpu_inst.shift_right ));
 sky130_fd_sc_hd__dfxtp_1 _2246_ (.CLK(clknet_4_2_0_clk),
    .D(_0099_),
    .Q(\cpu_inst.rotate ));
 sky130_fd_sc_hd__dfxtp_1 _2247_ (.CLK(clknet_4_2_0_clk),
    .D(_0100_),
    .Q(\cpu_inst.op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2248_ (.CLK(clknet_4_9_0_clk),
    .D(_0101_),
    .Q(\cpu_inst.op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2249_ (.CLK(clknet_4_3_0_clk),
    .D(_0102_),
    .Q(\cpu_inst.op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2250_ (.CLK(clknet_4_9_0_clk),
    .D(_0103_),
    .Q(\cpu_inst.op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2251_ (.CLK(clknet_4_9_0_clk),
    .D(_0104_),
    .Q(\cpu_inst.bit_ins ));
 sky130_fd_sc_hd__dfxtp_1 _2252_ (.CLK(clknet_4_8_0_clk),
    .D(_0105_),
    .Q(\cpu_inst.clv ));
 sky130_fd_sc_hd__dfxtp_1 _2253_ (.CLK(clknet_4_1_0_clk),
    .D(_0106_),
    .Q(\cpu_inst.sei ));
 sky130_fd_sc_hd__dfxtp_1 _2254_ (.CLK(clknet_4_0_0_clk),
    .D(_0107_),
    .Q(\cpu_inst.cli ));
 sky130_fd_sc_hd__dfxtp_1 _2255_ (.CLK(clknet_4_2_0_clk),
    .D(_0108_),
    .Q(\cpu_inst.sed ));
 sky130_fd_sc_hd__dfxtp_1 _2256_ (.CLK(clknet_4_3_0_clk),
    .D(_0109_),
    .Q(\cpu_inst.sec ));
 sky130_fd_sc_hd__dfxtp_1 _2257_ (.CLK(clknet_4_3_0_clk),
    .D(_0110_),
    .Q(\cpu_inst.clc ));
 sky130_fd_sc_hd__dfxtp_1 _2258_ (.CLK(clknet_4_3_0_clk),
    .D(_0111_),
    .Q(\cpu_inst.php ));
 sky130_fd_sc_hd__dfxtp_2 _2259_ (.CLK(clknet_4_1_0_clk),
    .D(_0112_),
    .Q(\cpu_inst.plp ));
 sky130_fd_sc_hd__dfxtp_1 _2260_ (.CLK(clknet_4_1_0_clk),
    .D(_0113_),
    .Q(\cpu_inst.cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2261_ (.CLK(clknet_4_8_0_clk),
    .D(_0114_),
    .Q(\cpu_inst.cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2262_ (.CLK(clknet_4_8_0_clk),
    .D(_0115_),
    .Q(\cpu_inst.cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2263_ (.CLK(clknet_4_12_0_clk),
    .D(_0116_),
    .Q(\cpu_inst.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2264_ (.CLK(clknet_4_12_0_clk),
    .D(_0117_),
    .Q(\cpu_inst.PC[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2265_ (.CLK(clknet_4_14_0_clk),
    .D(_0118_),
    .Q(\cpu_inst.PC[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2266_ (.CLK(clknet_4_14_0_clk),
    .D(_0119_),
    .Q(\cpu_inst.PC[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2267_ (.CLK(clknet_4_14_0_clk),
    .D(_0120_),
    .Q(\cpu_inst.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2268_ (.CLK(clknet_4_14_0_clk),
    .D(_0121_),
    .Q(\cpu_inst.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2269_ (.CLK(clknet_4_15_0_clk),
    .D(_0122_),
    .Q(\cpu_inst.PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2270_ (.CLK(clknet_4_15_0_clk),
    .D(_0123_),
    .Q(\cpu_inst.PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2271_ (.CLK(clknet_4_6_0_clk),
    .D(_0124_),
    .Q(\cpu_inst.PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2272_ (.CLK(clknet_4_6_0_clk),
    .D(_0125_),
    .Q(\cpu_inst.PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2273_ (.CLK(clknet_4_13_0_clk),
    .D(_0126_),
    .Q(\cpu_inst.PC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2274_ (.CLK(clknet_4_13_0_clk),
    .D(_0127_),
    .Q(\cpu_inst.PC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2275_ (.CLK(clknet_4_13_0_clk),
    .D(_0128_),
    .Q(\cpu_inst.PC[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2276_ (.CLK(clknet_4_12_0_clk),
    .D(_0129_),
    .Q(\cpu_inst.PC[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2277_ (.CLK(clknet_4_15_0_clk),
    .D(_0130_),
    .Q(\cpu_inst.PC[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2278_ (.CLK(clknet_4_13_0_clk),
    .D(_0131_),
    .Q(\cpu_inst.PC[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2279_ (.CLK(clknet_4_6_0_clk),
    .D(net3),
    .Q(\cpu_inst.NMI_1 ));
 sky130_fd_sc_hd__dfxtp_1 _2280_ (.CLK(clknet_4_6_0_clk),
    .D(net199),
    .Q(\cpu_inst.NMI_edge ));
 sky130_fd_sc_hd__dfxtp_1 _2281_ (.CLK(clknet_4_9_0_clk),
    .D(_0133_),
    .Q(\cpu_inst.AXYS[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2282_ (.CLK(clknet_4_8_0_clk),
    .D(_0134_),
    .Q(\cpu_inst.AXYS[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2283_ (.CLK(clknet_4_10_0_clk),
    .D(_0135_),
    .Q(\cpu_inst.AXYS[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2284_ (.CLK(clknet_4_10_0_clk),
    .D(_0136_),
    .Q(\cpu_inst.AXYS[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2285_ (.CLK(clknet_4_10_0_clk),
    .D(_0137_),
    .Q(\cpu_inst.AXYS[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2286_ (.CLK(clknet_4_11_0_clk),
    .D(_0138_),
    .Q(\cpu_inst.AXYS[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2287_ (.CLK(clknet_4_10_0_clk),
    .D(_0139_),
    .Q(\cpu_inst.AXYS[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2288_ (.CLK(clknet_4_10_0_clk),
    .D(_0140_),
    .Q(\cpu_inst.AXYS[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2289_ (.CLK(clknet_4_8_0_clk),
    .D(_0141_),
    .Q(\cpu_inst.AXYS[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2290_ (.CLK(clknet_4_8_0_clk),
    .D(_0142_),
    .Q(\cpu_inst.AXYS[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2291_ (.CLK(clknet_4_10_0_clk),
    .D(_0143_),
    .Q(\cpu_inst.AXYS[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2292_ (.CLK(clknet_4_10_0_clk),
    .D(_0144_),
    .Q(\cpu_inst.AXYS[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2293_ (.CLK(clknet_4_10_0_clk),
    .D(_0145_),
    .Q(\cpu_inst.AXYS[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2294_ (.CLK(clknet_4_11_0_clk),
    .D(_0146_),
    .Q(\cpu_inst.AXYS[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2295_ (.CLK(clknet_4_10_0_clk),
    .D(_0147_),
    .Q(\cpu_inst.AXYS[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2296_ (.CLK(clknet_4_10_0_clk),
    .D(_0148_),
    .Q(\cpu_inst.AXYS[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2297_ (.CLK(clknet_4_8_0_clk),
    .D(_0149_),
    .Q(\cpu_inst.AXYS[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2298_ (.CLK(clknet_4_8_0_clk),
    .D(_0150_),
    .Q(\cpu_inst.AXYS[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2299_ (.CLK(clknet_4_10_0_clk),
    .D(_0151_),
    .Q(\cpu_inst.AXYS[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2300_ (.CLK(clknet_4_10_0_clk),
    .D(_0152_),
    .Q(\cpu_inst.AXYS[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2301_ (.CLK(clknet_4_10_0_clk),
    .D(_0153_),
    .Q(\cpu_inst.AXYS[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2302_ (.CLK(clknet_4_11_0_clk),
    .D(_0154_),
    .Q(\cpu_inst.AXYS[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2303_ (.CLK(clknet_4_10_0_clk),
    .D(_0155_),
    .Q(\cpu_inst.AXYS[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2304_ (.CLK(clknet_4_10_0_clk),
    .D(_0156_),
    .Q(\cpu_inst.AXYS[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2305_ (.CLK(clknet_4_7_0_clk),
    .D(net142),
    .Q(\spi_sram_master_inst.data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2306_ (.CLK(clknet_4_7_0_clk),
    .D(_0158_),
    .Q(\spi_sram_master_inst.data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2307_ (.CLK(clknet_4_7_0_clk),
    .D(net150),
    .Q(\spi_sram_master_inst.data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2308_ (.CLK(clknet_4_6_0_clk),
    .D(_0160_),
    .Q(\spi_sram_master_inst.data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2309_ (.CLK(clknet_4_6_0_clk),
    .D(_0161_),
    .Q(\spi_sram_master_inst.data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2310_ (.CLK(clknet_4_6_0_clk),
    .D(_0162_),
    .Q(\spi_sram_master_inst.data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2311_ (.CLK(clknet_4_6_0_clk),
    .D(_0163_),
    .Q(\spi_sram_master_inst.data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2312_ (.CLK(clknet_4_7_0_clk),
    .D(net167),
    .Q(\spi_sram_master_inst.data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2313_ (.CLK(clknet_4_7_0_clk),
    .D(net127),
    .Q(\spi_sram_master_inst.data[33] ));
 sky130_fd_sc_hd__dfxtp_1 _2314_ (.CLK(clknet_4_7_0_clk),
    .D(_0166_),
    .Q(\spi_sram_master_inst.data[34] ));
 sky130_fd_sc_hd__dfxtp_1 _2315_ (.CLK(clknet_4_7_0_clk),
    .D(net139),
    .Q(\spi_sram_master_inst.data[35] ));
 sky130_fd_sc_hd__dfxtp_1 _2316_ (.CLK(clknet_4_7_0_clk),
    .D(_0168_),
    .Q(\spi_sram_master_inst.data[36] ));
 sky130_fd_sc_hd__dfxtp_1 _2317_ (.CLK(clknet_4_7_0_clk),
    .D(_0169_),
    .Q(\spi_sram_master_inst.data[37] ));
 sky130_fd_sc_hd__dfxtp_1 _2318_ (.CLK(clknet_4_7_0_clk),
    .D(net158),
    .Q(\spi_sram_master_inst.data[38] ));
 sky130_fd_sc_hd__dfxtp_1 _2319_ (.CLK(clknet_4_7_0_clk),
    .D(net125),
    .Q(\spi_sram_master_inst.data[39] ));
 sky130_fd_sc_hd__dfxtp_1 _2320_ (.CLK(clknet_4_4_0_clk),
    .D(_0172_),
    .Q(\spi_sram_master_inst.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2321_ (.CLK(clknet_4_4_0_clk),
    .D(_0173_),
    .Q(\spi_sram_master_inst.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2322_ (.CLK(clknet_4_4_0_clk),
    .D(_0174_),
    .Q(\spi_sram_master_inst.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2323_ (.CLK(clknet_4_5_0_clk),
    .D(_0175_),
    .Q(\spi_sram_master_inst.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2324_ (.CLK(clknet_4_11_0_clk),
    .D(_0176_),
    .Q(\cpu_inst.ALU.BI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2325_ (.CLK(net122),
    .D(\spi_sram_master_inst.data[39] ),
    .Q(\spi_sram_master_inst.dout ));
 sky130_fd_sc_hd__dfxtp_1 _2326_ (.CLK(net123),
    .D(\spi_sram_master_inst.cs_n_sm ),
    .Q(\spi_sram_master_inst.cs_n ));
 sky130_fd_sc_hd__dfxtp_1 _2327_ (.CLK(clknet_4_8_0_clk),
    .D(_0177_),
    .Q(\cpu_inst.AXYS[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2328_ (.CLK(clknet_4_8_0_clk),
    .D(_0178_),
    .Q(\cpu_inst.AXYS[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2329_ (.CLK(clknet_4_8_0_clk),
    .D(_0179_),
    .Q(\cpu_inst.AXYS[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2330_ (.CLK(clknet_4_10_0_clk),
    .D(_0180_),
    .Q(\cpu_inst.AXYS[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2331_ (.CLK(clknet_4_10_0_clk),
    .D(_0181_),
    .Q(\cpu_inst.AXYS[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2332_ (.CLK(clknet_4_11_0_clk),
    .D(_0182_),
    .Q(\cpu_inst.AXYS[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2333_ (.CLK(clknet_4_10_0_clk),
    .D(_0183_),
    .Q(\cpu_inst.AXYS[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2334_ (.CLK(clknet_4_10_0_clk),
    .D(_0184_),
    .Q(\cpu_inst.AXYS[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2335_ (.CLK(clknet_4_5_0_clk),
    .D(_0185_),
    .Q(\spi_sram_master_inst.counter_done ));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_121 (.HI(net121));
 sky130_fd_sc_hd__inv_2 _1087__1 (.A(clknet_4_5_0_clk),
    .Y(net122));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_119 (.HI(net119));
 sky130_fd_sc_hd__buf_2 _2357_ (.A(\spi_sram_master_inst.cs_n ),
    .X(uio_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _2358_ (.A(\spi_sram_master_inst.dout ),
    .X(uio_out[1]));
 sky130_fd_sc_hd__buf_2 _2359_ (.A(clknet_4_5_0_clk),
    .X(uio_out[3]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1198 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(ui_in[6]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[7]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(uio_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(_0274_),
    .X(net5));
 sky130_fd_sc_hd__buf_2 fanout6 (.A(_0274_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(_0902_),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 fanout8 (.A(net9),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 max_cap9 (.A(_0902_),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(_0985_),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(_0796_),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(_0795_),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net19),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(_0575_),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net23),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 fanout23 (.A(_0574_),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(_0365_),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(_0365_),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(_0807_),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net30),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(_0528_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net35),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net35),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(_0528_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net44),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net44),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net44),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net44),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(_0527_),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 wire45 (.A(_0808_),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(_0369_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(_0369_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 max_cap48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 wire49 (.A(_0803_),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(_0580_),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(_0685_),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(_0647_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net59),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net58),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(_0643_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(_0642_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(_0621_),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(_0579_),
    .X(net62));
 sky130_fd_sc_hd__buf_2 fanout63 (.A(_0579_),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_2 fanout65 (.A(_0572_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(_0537_),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(_0524_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 fanout70 (.A(_0523_),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(_0607_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(_0553_),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(_0553_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(_0534_),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(_0530_),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 fanout76 (.A(_0530_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(\cpu_inst.IRHOLD_valid ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(\cpu_inst.ADD[7] ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(\cpu_inst.ADD[6] ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(\cpu_inst.ADD[5] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(\cpu_inst.ADD[4] ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(\cpu_inst.ADD[3] ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(\cpu_inst.ADD[2] ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(\cpu_inst.ADD[1] ),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(\cpu_inst.ADD[0] ),
    .X(net85));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(\cpu_inst.state[3] ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(\cpu_inst.state[3] ),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(\cpu_inst.state[2] ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(\cpu_inst.state[2] ),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(\cpu_inst.state[1] ),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(\cpu_inst.state[0] ),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout93 (.A(\cpu_inst.state[0] ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 fanout94 (.A(\cpu_inst.DI[7] ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(\cpu_inst.DI[6] ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(\cpu_inst.DI[3] ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 fanout97 (.A(\cpu_inst.DI[2] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(\cpu_inst.DI[1] ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(\cpu_inst.DI[0] ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 fanout100 (.A(net1),
    .X(net100));
 sky130_fd_sc_hd__conb_1 tt_um_anders_tt_6502_101 (.LO(net101));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_12 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_6 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__inv_6 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\spi_sram_master_inst.data[39] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0171_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\spi_sram_master_inst.data[33] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0165_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\spi_sram_master_inst.counter[4] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\cpu_inst.IRHOLD[0] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\cpu_inst.AXYS[3][5] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\cpu_inst.AXYS[3][4] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\cpu_inst.AXYS[3][6] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\cpu_inst.AXYS[3][2] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\cpu_inst.AXYS[3][1] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\cpu_inst.IRHOLD[2] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\cpu_inst.AXYS[3][3] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\cpu_inst.dst_reg[0] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\spi_sram_master_inst.data[35] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0167_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\cpu_inst.IRHOLD[6] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\spi_sram_master_inst.data[24] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0157_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\cpu_inst.AXYS[0][1] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\cpu_inst.load_only ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\cpu_inst.AXYS[0][2] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\cpu_inst.src_reg[0] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\cpu_inst.AXYS[3][7] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\cpu_inst.AXYS[0][0] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\spi_sram_master_inst.data[26] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0159_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\cpu_inst.AXYS[0][6] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\spi_sram_master_inst.data[27] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\spi_sram_master_inst.data[36] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\cpu_inst.AXYS[0][4] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\cpu_inst.IRHOLD[5] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\cpu_inst.AXYS[2][1] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\spi_sram_master_inst.data[38] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0170_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\cpu_inst.dst_reg[1] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\spi_sram_master_inst.data[28] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\cpu_inst.AXYS[0][5] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\spi_sram_master_inst.data[34] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\cpu_inst.IRHOLD[3] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\cpu_inst.op[2] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\cpu_inst.IRHOLD[1] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\spi_sram_master_inst.data[31] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0164_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\cpu_inst.AXYS[0][3] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\spi_sram_master_inst.data[37] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\cpu_inst.res ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\spi_sram_master_inst.data[29] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\cpu_inst.index_y ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\cpu_inst.AXYS[2][4] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\cpu_inst.sed ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\cpu_inst.AXYS[1][3] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\cpu_inst.IRHOLD[7] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\cpu_inst.src_reg[1] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\cpu_inst.AXYS[1][4] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\cpu_inst.AXYS[2][7] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\cpu_inst.AXYS[2][5] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\cpu_inst.AXYS[1][5] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\cpu_inst.AXYS[1][1] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\cpu_inst.AXYS[0][7] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\cpu_inst.AXYS[3][0] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\cpu_inst.AXYS[2][2] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\cpu_inst.AXYS[2][6] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\cpu_inst.AXYS[2][3] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\spi_sram_master_inst.data[30] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\spi_sram_master_inst.data[25] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\cpu_inst.sec ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\cpu_inst.AXYS[1][7] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\cpu_inst.AXYS[2][0] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\cpu_inst.AXYS[1][6] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\spi_sram_master_inst.data[32] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\cpu_inst.sei ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\spi_sram_master_inst.counter[1] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0794_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\cpu_inst.NMI_1 ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0132_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\cpu_inst.ALU.AI7 ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\cpu_inst.inc ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\cpu_inst.ALU.BI7 ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\cpu_inst.ABL[0] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\cpu_inst.Z ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\cpu_inst.cond_code[0] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\spi_sram_master_inst.data[11] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\cpu_inst.ABL[1] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\cpu_inst.ABL[3] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\cpu_inst.ABL[2] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\spi_sram_master_inst.data[8] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\spi_sram_master_inst.data[17] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0031_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\spi_sram_master_inst.data[19] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0033_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\spi_sram_master_inst.data[9] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\spi_sram_master_inst.data[20] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\spi_sram_master_inst.data[15] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\spi_sram_master_inst.data[21] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\spi_sram_master_inst.data[22] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0036_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\cpu_inst.cond_code[2] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\spi_sram_master_inst.data[14] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\cpu_inst.store ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\spi_sram_master_inst.data[16] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\spi_sram_master_inst.data[12] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0026_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\cpu_inst.ABL[6] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\cpu_inst.AXYS[1][0] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\cpu_inst.ABL[5] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\spi_sram_master_inst.data[10] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0024_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\spi_sram_master_inst.data[13] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0027_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\spi_sram_master_inst.counter[0] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\spi_sram_master_inst.data[18] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\cpu_inst.bit_ins ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\cpu_inst.ABL[4] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\cpu_inst.N ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\cpu_inst.ABH[3] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\cpu_inst.IRHOLD[4] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\cpu_inst.cond_code[1] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\cpu_inst.shift ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\cpu_inst.V ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\cpu_inst.write_back ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\cpu_inst.clc ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\cpu_inst.ABH[4] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\cpu_inst.ABL[7] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\cpu_inst.ABH[1] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\cpu_inst.clv ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\cpu_inst.cld ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\cpu_inst.ABH[2] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\cpu_inst.ALU.HC ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\cpu_inst.cli ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\cpu_inst.D ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\cpu_inst.rotate ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\cpu_inst.PC[11] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\cpu_inst.AXYS[1][2] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\cpu_inst.PC[9] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\cpu_inst.PC[13] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\cpu_inst.load_reg ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\cpu_inst.adc_sbc ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\cpu_inst.PC[8] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\cpu_inst.PC[15] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\cpu_inst.PC[12] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\cpu_inst.PC[14] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\cpu_inst.PC[2] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\cpu_inst.PC[10] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\cpu_inst.PC[4] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\cpu_inst.op[0] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\spi_sram_master_inst.data[10] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\spi_sram_master_inst.data[14] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\spi_sram_master_inst.data[13] ),
    .X(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net54));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 assign uio_oe[0] = net119;
 assign uio_oe[1] = net120;
 assign uio_oe[2] = net101;
 assign uio_oe[3] = net121;
 assign uio_oe[4] = net102;
 assign uio_oe[5] = net103;
 assign uio_oe[6] = net104;
 assign uio_oe[7] = net105;
 assign uio_out[2] = net106;
 assign uio_out[4] = net107;
 assign uio_out[5] = net108;
 assign uio_out[6] = net109;
 assign uio_out[7] = net110;
 assign uo_out[0] = net111;
 assign uo_out[1] = net112;
 assign uo_out[2] = net113;
 assign uo_out[3] = net114;
 assign uo_out[4] = net115;
 assign uo_out[5] = net116;
 assign uo_out[6] = net117;
 assign uo_out[7] = net118;
endmodule
